`timescale 1ns / 1ps
    module rom (
    input clk,
    input en,
    input [12:0] addr,
    output reg [31:0] data
    );

    always @(posedge clk) begin
    if (en)
        case(addr)
			13'h0000: data <= 32'h00000000;	13'h0001: data <= 32'h0044A10B;	13'h0002: data <= 32'h00894204;	13'h0003: data <= 32'h00CDE2D4;	13'h0004: data <= 32'h0112836A;	13'h0005: data <= 32'h015723B1;	13'h0006: data <= 32'h019BC395;	13'h0007: data <= 32'h01E06302;	13'h0008: data <= 32'h022501E6;	13'h0009: data <= 32'h0269A02C;	13'h000A: data <= 32'h02AE3DC0;	13'h000B: data <= 32'h02F2DA8F;	13'h000C: data <= 32'h03377685;	13'h000D: data <= 32'h037C118E;	13'h000E: data <= 32'h03C0AB96;	13'h000F: data <= 32'h0405448B;	13'h0010: data <= 32'h0449DC58;	13'h0011: data <= 32'h048E72E9;	13'h0012: data <= 32'h04D3082A;	13'h0013: data <= 32'h05179C09;	13'h0014: data <= 32'h055C2E71;	13'h0015: data <= 32'h05A0BF4F;	13'h0016: data <= 32'h05E54E8E;	13'h0017: data <= 32'h0629DC1B;	13'h0018: data <= 32'h066E67E3;	13'h0019: data <= 32'h06B2F1D2;	13'h001A: data <= 32'h06F779D3;	13'h001B: data <= 32'h073BFFD4;	13'h001C: data <= 32'h078083C0;	13'h001D: data <= 32'h07C50585;	13'h001E: data <= 32'h0809850D;	13'h001F: data <= 32'h084E0246;	13'h0020: data <= 32'h08927D1C;	13'h0021: data <= 32'h08D6F57B;	13'h0022: data <= 32'h091B6B50;	13'h0023: data <= 32'h095FDE86;	13'h0024: data <= 32'h09A44F0B;	13'h0025: data <= 32'h09E8BCC9;	13'h0026: data <= 32'h0A2D27AF;	13'h0027: data <= 32'h0A718FA8;	13'h0028: data <= 32'h0AB5F4A0;	13'h0029: data <= 32'h0AFA5684;	13'h002A: data <= 32'h0B3EB53F;	13'h002B: data <= 32'h0B8310C0;	13'h002C: data <= 32'h0BC768F1;	13'h002D: data <= 32'h0C0BBDBF;	13'h002E: data <= 32'h0C500F17;	13'h002F: data <= 32'h0C945CE5;	13'h0030: data <= 32'h0CD8A715;	13'h0031: data <= 32'h0D1CED93;	13'h0032: data <= 32'h0D61304D;	13'h0033: data <= 32'h0DA56F2E;	13'h0034: data <= 32'h0DE9AA23;	13'h0035: data <= 32'h0E2DE117;	13'h0036: data <= 32'h0E7213F8;	13'h0037: data <= 32'h0EB642B3;	13'h0038: data <= 32'h0EFA6D32;	13'h0039: data <= 32'h0F3E9363;	13'h003A: data <= 32'h0F82B532;	13'h003B: data <= 32'h0FC6D28C;	13'h003C: data <= 32'h100AEB5D;	13'h003D: data <= 32'h104EFF91;	13'h003E: data <= 32'h10930F15;	13'h003F: data <= 32'h10D719D5;	13'h0040: data <= 32'h111B1FBE;	13'h0041: data <= 32'h115F20BC;	13'h0042: data <= 32'h11A31CBB;	13'h0043: data <= 32'h11E713A9;	13'h0044: data <= 32'h122B0571;	13'h0045: data <= 32'h126EF200;	13'h0046: data <= 32'h12B2D942;	13'h0047: data <= 32'h12F6BB25;	13'h0048: data <= 32'h133A9793;	13'h0049: data <= 32'h137E6E7B;	13'h004A: data <= 32'h13C23FC8;	13'h004B: data <= 32'h14060B67;	13'h004C: data <= 32'h1449D144;	13'h004D: data <= 32'h148D914D;	13'h004E: data <= 32'h14D14B6C;	13'h004F: data <= 32'h1514FF90;	13'h0050: data <= 32'h1558ADA4;	13'h0051: data <= 32'h159C5595;	13'h0052: data <= 32'h15DFF750;	13'h0053: data <= 32'h162392C1;	13'h0054: data <= 32'h166727D4;	13'h0055: data <= 32'h16AAB677;	13'h0056: data <= 32'h16EE3E96;	13'h0057: data <= 32'h1731C01E;	13'h0058: data <= 32'h17753AFA;	13'h0059: data <= 32'h17B8AF18;	13'h005A: data <= 32'h17FC1C64;	13'h005B: data <= 32'h183F82CC;	13'h005C: data <= 32'h1882E23A;	13'h005D: data <= 32'h18C63A9D;	13'h005E: data <= 32'h19098BE1;	13'h005F: data <= 32'h194CD5F2;	13'h0060: data <= 32'h199018BD;	13'h0061: data <= 32'h19D3542F;	13'h0062: data <= 32'h1A168834;	13'h0063: data <= 32'h1A59B4B9;	13'h0064: data <= 32'h1A9CD9AC;	13'h0065: data <= 32'h1ADFF6F7;	13'h0066: data <= 32'h1B230C89;	13'h0067: data <= 32'h1B661A4E;	13'h0068: data <= 32'h1BA92032;	13'h0069: data <= 32'h1BEC1E23;	13'h006A: data <= 32'h1C2F140D;	13'h006B: data <= 32'h1C7201DD;	13'h006C: data <= 32'h1CB4E77F;	13'h006D: data <= 32'h1CF7C4E1;	13'h006E: data <= 32'h1D3A99EF;	13'h006F: data <= 32'h1D7D6696;	13'h0070: data <= 32'h1DC02AC2;	13'h0071: data <= 32'h1E02E662;	13'h0072: data <= 32'h1E459960;	13'h0073: data <= 32'h1E8843AB;	13'h0074: data <= 32'h1ECAE52F;	13'h0075: data <= 32'h1F0D7DD8;	13'h0076: data <= 32'h1F500D95;	13'h0077: data <= 32'h1F929451;	13'h0078: data <= 32'h1FD511F9;	13'h0079: data <= 32'h2017867B;	13'h007A: data <= 32'h2059F1C3;	13'h007B: data <= 32'h209C53BF;	13'h007C: data <= 32'h20DEAC5A;	13'h007D: data <= 32'h2120FB82;	13'h007E: data <= 32'h21634125;	13'h007F: data <= 32'h21A57D2E;	13'h0080: data <= 32'h21E7AF8B;	13'h0081: data <= 32'h2229D829;	13'h0082: data <= 32'h226BF6F5;	13'h0083: data <= 32'h22AE0BDB;	13'h0084: data <= 32'h22F016C9;	13'h0085: data <= 32'h233217AD;	13'h0086: data <= 32'h23740E72;	13'h0087: data <= 32'h23B5FB05;	13'h0088: data <= 32'h23F7DD55;	13'h0089: data <= 32'h2439B54E;	13'h008A: data <= 32'h247B82DD;	13'h008B: data <= 32'h24BD45EF;	13'h008C: data <= 32'h24FEFE71;	13'h008D: data <= 32'h2540AC50;	13'h008E: data <= 32'h25824F7A;	13'h008F: data <= 32'h25C3E7DC;	13'h0090: data <= 32'h26057562;	13'h0091: data <= 32'h2646F7FB;	13'h0092: data <= 32'h26886F92;	13'h0093: data <= 32'h26C9DC16;	13'h0094: data <= 32'h270B3D72;	13'h0095: data <= 32'h274C9396;	13'h0096: data <= 32'h278DDE6E;	13'h0097: data <= 32'h27CF1DE6;	13'h0098: data <= 32'h281051ED;	13'h0099: data <= 32'h28517A6F;	13'h009A: data <= 32'h2892975B;	13'h009B: data <= 32'h28D3A89C;	13'h009C: data <= 32'h2914AE21;	13'h009D: data <= 32'h2955A7D7;	13'h009E: data <= 32'h299695AA;	13'h009F: data <= 32'h29D7778A;	13'h00A0: data <= 32'h2A184D61;	13'h00A1: data <= 32'h2A59171F;	13'h00A2: data <= 32'h2A99D4B1;	13'h00A3: data <= 32'h2ADA8603;	13'h00A4: data <= 32'h2B1B2B04;	13'h00A5: data <= 32'h2B5BC3A0;	13'h00A6: data <= 32'h2B9C4FC5;	13'h00A7: data <= 32'h2BDCCF61;	13'h00A8: data <= 32'h2C1D4261;	13'h00A9: data <= 32'h2C5DA8B3;	13'h00AA: data <= 32'h2C9E0243;	13'h00AB: data <= 32'h2CDE4F00;	13'h00AC: data <= 32'h2D1E8ED7;	13'h00AD: data <= 32'h2D5EC1B5;	13'h00AE: data <= 32'h2D9EE789;	13'h00AF: data <= 32'h2DDF003F;	13'h00B0: data <= 32'h2E1F0BC5;	13'h00B1: data <= 32'h2E5F0A09;	13'h00B2: data <= 32'h2E9EFAF9;	13'h00B3: data <= 32'h2EDEDE81;	13'h00B4: data <= 32'h2F1EB490;	13'h00B5: data <= 32'h2F5E7D14;	13'h00B6: data <= 32'h2F9E37F9;	13'h00B7: data <= 32'h2FDDE52E;	13'h00B8: data <= 32'h301D84A1;	13'h00B9: data <= 32'h305D163E;	13'h00BA: data <= 32'h309C99F5;	13'h00BB: data <= 32'h30DC0FB1;	13'h00BC: data <= 32'h311B7762;	13'h00BD: data <= 32'h315AD0F5;	13'h00BE: data <= 32'h319A1C58;	13'h00BF: data <= 32'h31D95979;	13'h00C0: data <= 32'h32188845;	13'h00C1: data <= 32'h3257A8AA;	13'h00C2: data <= 32'h3296BA97;	13'h00C3: data <= 32'h32D5BDF8;	13'h00C4: data <= 32'h3314B2BC;	13'h00C5: data <= 32'h335398D2;	13'h00C6: data <= 32'h33927025;	13'h00C7: data <= 32'h33D138A6;	13'h00C8: data <= 32'h340FF241;	13'h00C9: data <= 32'h344E9CE5;	13'h00CA: data <= 32'h348D387F;	13'h00CB: data <= 32'h34CBC4FE;	13'h00CC: data <= 32'h350A424F;	13'h00CD: data <= 32'h3548B061;	13'h00CE: data <= 32'h35870F22;	13'h00CF: data <= 32'h35C55E80;	13'h00D0: data <= 32'h36039E68;	13'h00D1: data <= 32'h3641CEC9;	13'h00D2: data <= 32'h367FEF91;	13'h00D3: data <= 32'h36BE00AF;	13'h00D4: data <= 32'h36FC0210;	13'h00D5: data <= 32'h3739F3A2;	13'h00D6: data <= 32'h3777D554;	13'h00D7: data <= 32'h37B5A714;	13'h00D8: data <= 32'h37F368D0;	13'h00D9: data <= 32'h38311A77;	13'h00DA: data <= 32'h386EBBF6;	13'h00DB: data <= 32'h38AC4D3C;	13'h00DC: data <= 32'h38E9CE38;	13'h00DD: data <= 32'h39273ED7;	13'h00DE: data <= 32'h39649F08;	13'h00DF: data <= 32'h39A1EEB9;	13'h00E0: data <= 32'h39DF2DD9;	13'h00E1: data <= 32'h3A1C5C56;	13'h00E2: data <= 32'h3A597A1E;	13'h00E3: data <= 32'h3A968720;	13'h00E4: data <= 32'h3AD3834B;	13'h00E5: data <= 32'h3B106E8C;	13'h00E6: data <= 32'h3B4D48D3;	13'h00E7: data <= 32'h3B8A120D;	13'h00E8: data <= 32'h3BC6CA2A;	13'h00E9: data <= 32'h3C037117;	13'h00EA: data <= 32'h3C4006C4;	13'h00EB: data <= 32'h3C7C8B1F;	13'h00EC: data <= 32'h3CB8FE17;	13'h00ED: data <= 32'h3CF55F9A;	13'h00EE: data <= 32'h3D31AF97;	13'h00EF: data <= 32'h3D6DEDFC;	13'h00F0: data <= 32'h3DAA1AB9;	13'h00F1: data <= 32'h3DE635BB;	13'h00F2: data <= 32'h3E223EF2;	13'h00F3: data <= 32'h3E5E364C;	13'h00F4: data <= 32'h3E9A1BB9;	13'h00F5: data <= 32'h3ED5EF27;	13'h00F6: data <= 32'h3F11B084;	13'h00F7: data <= 32'h3F4D5FC0;	13'h00F8: data <= 32'h3F88FCC9;	13'h00F9: data <= 32'h3FC4878E;	13'h00FA: data <= 32'h3FFFFFFF;	13'h00FB: data <= 32'h403B660A;	13'h00FC: data <= 32'h4076B99D;	13'h00FD: data <= 32'h40B1FAA9;	13'h00FE: data <= 32'h40ED291B;	13'h00FF: data <= 32'h412844E3;	13'h0100: data <= 32'h41634DF1;	13'h0101: data <= 32'h419E4432;	13'h0102: data <= 32'h41D92796;	13'h0103: data <= 32'h4213F80C;	13'h0104: data <= 32'h424EB583;	13'h0105: data <= 32'h42895FEA;	13'h0106: data <= 32'h42C3F731;	13'h0107: data <= 32'h42FE7B46;	13'h0108: data <= 32'h4338EC19;	13'h0109: data <= 32'h43734999;	13'h010A: data <= 32'h43AD93B5;	13'h010B: data <= 32'h43E7CA5C;	13'h010C: data <= 32'h4421ED7E;	13'h010D: data <= 32'h445BFD0A;	13'h010E: data <= 32'h4495F8EF;	13'h010F: data <= 32'h44CFE11D;	13'h0110: data <= 32'h4509B583;	13'h0111: data <= 32'h4543760F;	13'h0112: data <= 32'h457D22B3;	13'h0113: data <= 32'h45B6BB5D;	13'h0114: data <= 32'h45F03FFC;	13'h0115: data <= 32'h4629B080;	13'h0116: data <= 32'h46630CD9;	13'h0117: data <= 32'h469C54F6;	13'h0118: data <= 32'h46D588C6;	13'h0119: data <= 32'h470EA839;	13'h011A: data <= 32'h4747B33F;	13'h011B: data <= 32'h4780A9C8;	13'h011C: data <= 32'h47B98BC2;	13'h011D: data <= 32'h47F2591E;	13'h011E: data <= 32'h482B11CB;	13'h011F: data <= 32'h4863B5B9;	13'h0120: data <= 32'h489C44D7;	13'h0121: data <= 32'h48D4BF16;	13'h0122: data <= 32'h490D2465;	13'h0123: data <= 32'h494574B4;	13'h0124: data <= 32'h497DAFF3;	13'h0125: data <= 32'h49B5D611;	13'h0126: data <= 32'h49EDE6FF;	13'h0127: data <= 32'h4A25E2AC;	13'h0128: data <= 32'h4A5DC908;	13'h0129: data <= 32'h4A959A04;	13'h012A: data <= 32'h4ACD558E;	13'h012B: data <= 32'h4B04FB98;	13'h012C: data <= 32'h4B3C8C11;	13'h012D: data <= 32'h4B7406E9;	13'h012E: data <= 32'h4BAB6C10;	13'h012F: data <= 32'h4BE2BB76;	13'h0130: data <= 32'h4C19F50B;	13'h0131: data <= 32'h4C5118C0;	13'h0132: data <= 32'h4C882685;	13'h0133: data <= 32'h4CBF1E4A;	13'h0134: data <= 32'h4CF5FFFE;	13'h0135: data <= 32'h4D2CCB93;	13'h0136: data <= 32'h4D6380F8;	13'h0137: data <= 32'h4D9A201D;	13'h0138: data <= 32'h4DD0A8F4;	13'h0139: data <= 32'h4E071B6D;	13'h013A: data <= 32'h4E3D7776;	13'h013B: data <= 32'h4E73BD02;	13'h013C: data <= 32'h4EA9EC01;	13'h013D: data <= 32'h4EE00462;	13'h013E: data <= 32'h4F160617;	13'h013F: data <= 32'h4F4BF10F;	13'h0140: data <= 32'h4F81C53C;	13'h0141: data <= 32'h4FB7828E;	13'h0142: data <= 32'h4FED28F5;	13'h0143: data <= 32'h5022B862;	13'h0144: data <= 32'h505830C5;	13'h0145: data <= 32'h508D9210;	13'h0146: data <= 32'h50C2DC33;	13'h0147: data <= 32'h50F80F1E;	13'h0148: data <= 32'h512D2AC2;	13'h0149: data <= 32'h51622F11;	13'h014A: data <= 32'h51971BFA;	13'h014B: data <= 32'h51CBF16E;	13'h014C: data <= 32'h5200AF5F;	13'h014D: data <= 32'h523555BD;	13'h014E: data <= 32'h5269E47A;	13'h014F: data <= 32'h529E5B85;	13'h0150: data <= 32'h52D2BAD0;	13'h0151: data <= 32'h5307024B;	13'h0152: data <= 32'h533B31E9;	13'h0153: data <= 32'h536F4999;	13'h0154: data <= 32'h53A3494D;	13'h0155: data <= 32'h53D730F6;	13'h0156: data <= 32'h540B0085;	13'h0157: data <= 32'h543EB7EB;	13'h0158: data <= 32'h54725719;	13'h0159: data <= 32'h54A5DE00;	13'h015A: data <= 32'h54D94C92;	13'h015B: data <= 32'h550CA2BF;	13'h015C: data <= 32'h553FE07A;	13'h015D: data <= 32'h557305B2;	13'h015E: data <= 32'h55A6125A;	13'h015F: data <= 32'h55D90663;	13'h0160: data <= 32'h560BE1BF;	13'h0161: data <= 32'h563EA45D;	13'h0162: data <= 32'h56714E31;	13'h0163: data <= 32'h56A3DF2B;	13'h0164: data <= 32'h56D6573E;	13'h0165: data <= 32'h5708B659;	13'h0166: data <= 32'h573AFC6F;	13'h0167: data <= 32'h576D2972;	13'h0168: data <= 32'h579F3D53;	13'h0169: data <= 32'h57D13804;	13'h016A: data <= 32'h58031975;	13'h016B: data <= 32'h5834E19A;	13'h016C: data <= 32'h58669063;	13'h016D: data <= 32'h589825C3;	13'h016E: data <= 32'h58C9A1AA;	13'h016F: data <= 32'h58FB040C;	13'h0170: data <= 32'h592C4CD9;	13'h0171: data <= 32'h595D7C04;	13'h0172: data <= 32'h598E917E;	13'h0173: data <= 32'h59BF8D39;	13'h0174: data <= 32'h59F06F27;	13'h0175: data <= 32'h5A21373B;	13'h0176: data <= 32'h5A51E565;	13'h0177: data <= 32'h5A827999;	13'h0178: data <= 32'h5AB2F3C7;	13'h0179: data <= 32'h5AE353E3;	13'h017A: data <= 32'h5B1399DF;	13'h017B: data <= 32'h5B43C5AB;	13'h017C: data <= 32'h5B73D73B;	13'h017D: data <= 32'h5BA3CE81;	13'h017E: data <= 32'h5BD3AB6F;	13'h017F: data <= 32'h5C036DF7;	13'h0180: data <= 32'h5C33160B;	13'h0181: data <= 32'h5C62A39E;	13'h0182: data <= 32'h5C9216A3;	13'h0183: data <= 32'h5CC16F0A;	13'h0184: data <= 32'h5CF0ACC8;	13'h0185: data <= 32'h5D1FCFCE;	13'h0186: data <= 32'h5D4ED80E;	13'h0187: data <= 32'h5D7DC57C;	13'h0188: data <= 32'h5DAC9809;	13'h0189: data <= 32'h5DDB4FA9;	13'h018A: data <= 32'h5E09EC4D;	13'h018B: data <= 32'h5E386DE9;	13'h018C: data <= 32'h5E66D46E;	13'h018D: data <= 32'h5E951FD1;	13'h018E: data <= 32'h5EC35003;	13'h018F: data <= 32'h5EF164F7;	13'h0190: data <= 32'h5F1F5EA0;	13'h0191: data <= 32'h5F4D3CF0;	13'h0192: data <= 32'h5F7AFFDB;	13'h0193: data <= 32'h5FA8A753;	13'h0194: data <= 32'h5FD6334C;	13'h0195: data <= 32'h6003A3B7;	13'h0196: data <= 32'h6030F888;	13'h0197: data <= 32'h605E31B3;	13'h0198: data <= 32'h608B4F29;	13'h0199: data <= 32'h60B850DF;	13'h019A: data <= 32'h60E536C6;	13'h019B: data <= 32'h611200D3;	13'h019C: data <= 32'h613EAEF8;	13'h019D: data <= 32'h616B4129;	13'h019E: data <= 32'h6197B758;	13'h019F: data <= 32'h61C41179;	13'h01A0: data <= 32'h61F04F7F;	13'h01A1: data <= 32'h621C715D;	13'h01A2: data <= 32'h62487707;	13'h01A3: data <= 32'h62746071;	13'h01A4: data <= 32'h62A02D8C;	13'h01A5: data <= 32'h62CBDE4E;	13'h01A6: data <= 32'h62F772A8;	13'h01A7: data <= 32'h6322EA90;	13'h01A8: data <= 32'h634E45F8;	13'h01A9: data <= 32'h637984D3;	13'h01AA: data <= 32'h63A4A716;	13'h01AB: data <= 32'h63CFACB4;	13'h01AC: data <= 32'h63FA95A0;	13'h01AD: data <= 32'h642561CF;	13'h01AE: data <= 32'h64501133;	13'h01AF: data <= 32'h647AA3C2;	13'h01B0: data <= 32'h64A5196D;	13'h01B1: data <= 32'h64CF722A;	13'h01B2: data <= 32'h64F9ADEC;	13'h01B3: data <= 32'h6523CCA7;	13'h01B4: data <= 32'h654DCE4F;	13'h01B5: data <= 32'h6577B2D7;	13'h01B6: data <= 32'h65A17A34;	13'h01B7: data <= 32'h65CB245A;	13'h01B8: data <= 32'h65F4B13D;	13'h01B9: data <= 32'h661E20D0;	13'h01BA: data <= 32'h66477308;	13'h01BB: data <= 32'h6670A7D9;	13'h01BC: data <= 32'h6699BF37;	13'h01BD: data <= 32'h66C2B917;	13'h01BE: data <= 32'h66EB956C;	13'h01BF: data <= 32'h6714542B;	13'h01C0: data <= 32'h673CF548;	13'h01C1: data <= 32'h676578B7;	13'h01C2: data <= 32'h678DDE6D;	13'h01C3: data <= 32'h67B6265E;	13'h01C4: data <= 32'h67DE507F;	13'h01C5: data <= 32'h68065CC4;	13'h01C6: data <= 32'h682E4B21;	13'h01C7: data <= 32'h68561B8B;	13'h01C8: data <= 32'h687DCDF7;	13'h01C9: data <= 32'h68A56259;	13'h01CA: data <= 32'h68CCD8A5;	13'h01CB: data <= 32'h68F430D2;	13'h01CC: data <= 32'h691B6AD2;	13'h01CD: data <= 32'h6942869B;	13'h01CE: data <= 32'h69698422;	13'h01CF: data <= 32'h6990635B;	13'h01D0: data <= 32'h69B7243B;	13'h01D1: data <= 32'h69DDC6B8;	13'h01D2: data <= 32'h6A044AC5;	13'h01D3: data <= 32'h6A2AB058;	13'h01D4: data <= 32'h6A50F766;	13'h01D5: data <= 32'h6A771FE4;	13'h01D6: data <= 32'h6A9D29C7;	13'h01D7: data <= 32'h6AC31504;	13'h01D8: data <= 32'h6AE8E190;	13'h01D9: data <= 32'h6B0E8F60;	13'h01DA: data <= 32'h6B341E69;	13'h01DB: data <= 32'h6B598EA1;	13'h01DC: data <= 32'h6B7EDFFD;	13'h01DD: data <= 32'h6BA41272;	13'h01DE: data <= 32'h6BC925F5;	13'h01DF: data <= 32'h6BEE1A7C;	13'h01E0: data <= 32'h6C12EFFC;	13'h01E1: data <= 32'h6C37A66B;	13'h01E2: data <= 32'h6C5C3DBD;	13'h01E3: data <= 32'h6C80B5E9;	13'h01E4: data <= 32'h6CA50EE4;	13'h01E5: data <= 32'h6CC948A3;	13'h01E6: data <= 32'h6CED631D;	13'h01E7: data <= 32'h6D115E46;	13'h01E8: data <= 32'h6D353A15;	13'h01E9: data <= 32'h6D58F67E;	13'h01EA: data <= 32'h6D7C9378;	13'h01EB: data <= 32'h6DA010F9;	13'h01EC: data <= 32'h6DC36EF7;	13'h01ED: data <= 32'h6DE6AD66;	13'h01EE: data <= 32'h6E09CC3D;	13'h01EF: data <= 32'h6E2CCB73;	13'h01F0: data <= 32'h6E4FAAFC;	13'h01F1: data <= 32'h6E726ACF;	13'h01F2: data <= 32'h6E950AE2;	13'h01F3: data <= 32'h6EB78B2B;	13'h01F4: data <= 32'h6ED9EBA0;	13'h01F5: data <= 32'h6EFC2C37;	13'h01F6: data <= 32'h6F1E4CE6;	13'h01F7: data <= 32'h6F404DA4;	13'h01F8: data <= 32'h6F622E67;	13'h01F9: data <= 32'h6F83EF24;	13'h01FA: data <= 32'h6FA58FD3;	13'h01FB: data <= 32'h6FC71069;	13'h01FC: data <= 32'h6FE870DD;	13'h01FD: data <= 32'h7009B125;	13'h01FE: data <= 32'h702AD139;	13'h01FF: data <= 32'h704BD10D;	13'h0200: data <= 32'h706CB09A;	13'h0201: data <= 32'h708D6FD4;	13'h0202: data <= 32'h70AE0EB4;	13'h0203: data <= 32'h70CE8D2F;	13'h0204: data <= 32'h70EEEB3C;	13'h0205: data <= 32'h710F28D2;	13'h0206: data <= 32'h712F45E8;	13'h0207: data <= 32'h714F4274;	13'h0208: data <= 32'h716F1E6E;	13'h0209: data <= 32'h718ED9CB;	13'h020A: data <= 32'h71AE7484;	13'h020B: data <= 32'h71CDEE8E;	13'h020C: data <= 32'h71ED47E1;	13'h020D: data <= 32'h720C8074;	13'h020E: data <= 32'h722B983D;	13'h020F: data <= 32'h724A8F35;	13'h0210: data <= 32'h72696551;	13'h0211: data <= 32'h72881A89;	13'h0212: data <= 32'h72A6AED5;	13'h0213: data <= 32'h72C5222B;	13'h0214: data <= 32'h72E37483;	13'h0215: data <= 32'h7301A5D4;	13'h0216: data <= 32'h731FB615;	13'h0217: data <= 32'h733DA53E;	13'h0218: data <= 32'h735B7346;	13'h0219: data <= 32'h73792025;	13'h021A: data <= 32'h7396ABD1;	13'h021B: data <= 32'h73B41643;	13'h021C: data <= 32'h73D15F72;	13'h021D: data <= 32'h73EE8756;	13'h021E: data <= 32'h740B8DE5;	13'h021F: data <= 32'h74287319;	13'h0220: data <= 32'h744536E8;	13'h0221: data <= 32'h7461D94B;	13'h0222: data <= 32'h747E5A39;	13'h0223: data <= 32'h749AB9A9;	13'h0224: data <= 32'h74B6F794;	13'h0225: data <= 32'h74D313F2;	13'h0226: data <= 32'h74EF0EBB;	13'h0227: data <= 32'h750AE7E5;	13'h0228: data <= 32'h75269F6B;	13'h0229: data <= 32'h75423543;	13'h022A: data <= 32'h755DA965;	13'h022B: data <= 32'h7578FBCA;	13'h022C: data <= 32'h75942C6A;	13'h022D: data <= 32'h75AF3B3D;	13'h022E: data <= 32'h75CA283B;	13'h022F: data <= 32'h75E4F35D;	13'h0230: data <= 32'h75FF9C9A;	13'h0231: data <= 32'h761A23EC;	13'h0232: data <= 32'h7634894A;	13'h0233: data <= 32'h764ECCAD;	13'h0234: data <= 32'h7668EE0D;	13'h0235: data <= 32'h7682ED64;	13'h0236: data <= 32'h769CCAA8;	13'h0237: data <= 32'h76B685D4;	13'h0238: data <= 32'h76D01EDF;	13'h0239: data <= 32'h76E995C2;	13'h023A: data <= 32'h7702EA76;	13'h023B: data <= 32'h771C1CF4;	13'h023C: data <= 32'h77352D34;	13'h023D: data <= 32'h774E1B2F;	13'h023E: data <= 32'h7766E6DF;	13'h023F: data <= 32'h777F903B;	13'h0240: data <= 32'h7798173C;	13'h0241: data <= 32'h77B07BDD;	13'h0242: data <= 32'h77C8BE15;	13'h0243: data <= 32'h77E0DDDE;	13'h0244: data <= 32'h77F8DB31;	13'h0245: data <= 32'h7810B606;	13'h0246: data <= 32'h78286E58;	13'h0247: data <= 32'h7840041E;	13'h0248: data <= 32'h78577754;	13'h0249: data <= 32'h786EC7F1;	13'h024A: data <= 32'h7885F5EE;	13'h024B: data <= 32'h789D0147;	13'h024C: data <= 32'h78B3E9F3;	13'h024D: data <= 32'h78CAAFEC;	13'h024E: data <= 32'h78E1532B;	13'h024F: data <= 32'h78F7D3AB;	13'h0250: data <= 32'h790E3164;	13'h0251: data <= 32'h79246C50;	13'h0252: data <= 32'h793A846A;	13'h0253: data <= 32'h795079A9;	13'h0254: data <= 32'h79664C09;	13'h0255: data <= 32'h797BFB82;	13'h0256: data <= 32'h7991880F;	13'h0257: data <= 32'h79A6F1AA;	13'h0258: data <= 32'h79BC384C;	13'h0259: data <= 32'h79D15BEE;	13'h025A: data <= 32'h79E65C8C;	13'h025B: data <= 32'h79FB3A1F;	13'h025C: data <= 32'h7A0FF4A1;	13'h025D: data <= 32'h7A248C0C;	13'h025E: data <= 32'h7A39005A;	13'h025F: data <= 32'h7A4D5186;	13'h0260: data <= 32'h7A617F89;	13'h0261: data <= 32'h7A758A5D;	13'h0262: data <= 32'h7A8971FD;	13'h0263: data <= 32'h7A9D3664;	13'h0264: data <= 32'h7AB0D78B;	13'h0265: data <= 32'h7AC4556C;	13'h0266: data <= 32'h7AD7B003;	13'h0267: data <= 32'h7AEAE74A;	13'h0268: data <= 32'h7AFDFB3A;	13'h0269: data <= 32'h7B10EBD0;	13'h026A: data <= 32'h7B23B904;	13'h026B: data <= 32'h7B3662D2;	13'h026C: data <= 32'h7B48E935;	13'h026D: data <= 32'h7B5B4C27;	13'h026E: data <= 32'h7B6D8BA2;	13'h026F: data <= 32'h7B7FA7A3;	13'h0270: data <= 32'h7B91A022;	13'h0271: data <= 32'h7BA3751C;	13'h0272: data <= 32'h7BB5268A;	13'h0273: data <= 32'h7BC6B469;	13'h0274: data <= 32'h7BD81EB3;	13'h0275: data <= 32'h7BE96562;	13'h0276: data <= 32'h7BFA8873;	13'h0277: data <= 32'h7C0B87DF;	13'h0278: data <= 32'h7C1C63A3;	13'h0279: data <= 32'h7C2D1BB9;	13'h027A: data <= 32'h7C3DB01C;	13'h027B: data <= 32'h7C4E20C9;	13'h027C: data <= 32'h7C5E6DB9;	13'h027D: data <= 32'h7C6E96E8;	13'h027E: data <= 32'h7C7E9C53;	13'h027F: data <= 32'h7C8E7DF3;	13'h0280: data <= 32'h7C9E3BC4;	13'h0281: data <= 32'h7CADD5C3;	13'h0282: data <= 32'h7CBD4BEA;	13'h0283: data <= 32'h7CCC9E36;	13'h0284: data <= 32'h7CDBCCA0;	13'h0285: data <= 32'h7CEAD727;	13'h0286: data <= 32'h7CF9BDC4;	13'h0287: data <= 32'h7D088073;	13'h0288: data <= 32'h7D171F32;	13'h0289: data <= 32'h7D2599FA;	13'h028A: data <= 32'h7D33F0C8;	13'h028B: data <= 32'h7D422399;	13'h028C: data <= 32'h7D503267;	13'h028D: data <= 32'h7D5E1D2F;	13'h028E: data <= 32'h7D6BE3ED;	13'h028F: data <= 32'h7D79869D;	13'h0290: data <= 32'h7D87053A;	13'h0291: data <= 32'h7D945FC2;	13'h0292: data <= 32'h7DA19630;	13'h0293: data <= 32'h7DAEA880;	13'h0294: data <= 32'h7DBB96AF;	13'h0295: data <= 32'h7DC860B9;	13'h0296: data <= 32'h7DD5069A;	13'h0297: data <= 32'h7DE1884F;	13'h0298: data <= 32'h7DEDE5D4;	13'h0299: data <= 32'h7DFA1F25;	13'h029A: data <= 32'h7E06343F;	13'h029B: data <= 32'h7E12251F;	13'h029C: data <= 32'h7E1DF1C1;	13'h029D: data <= 32'h7E299A21;	13'h029E: data <= 32'h7E351E3D;	13'h029F: data <= 32'h7E407E11;	13'h02A0: data <= 32'h7E4BB999;	13'h02A1: data <= 32'h7E56D0D3;	13'h02A2: data <= 32'h7E61C3BC;	13'h02A3: data <= 32'h7E6C924F;	13'h02A4: data <= 32'h7E773C8B;	13'h02A5: data <= 32'h7E81C26B;	13'h02A6: data <= 32'h7E8C23EE;	13'h02A7: data <= 32'h7E96610F;	13'h02A8: data <= 32'h7EA079CD;	13'h02A9: data <= 32'h7EAA6E24;	13'h02AA: data <= 32'h7EB43E11;	13'h02AB: data <= 32'h7EBDE991;	13'h02AC: data <= 32'h7EC770A2;	13'h02AD: data <= 32'h7ED0D341;	13'h02AE: data <= 32'h7EDA116B;	13'h02AF: data <= 32'h7EE32B1E;	13'h02B0: data <= 32'h7EEC2057;	13'h02B1: data <= 32'h7EF4F113;	13'h02B2: data <= 32'h7EFD9D51;	13'h02B3: data <= 32'h7F06250C;	13'h02B4: data <= 32'h7F0E8843;	13'h02B5: data <= 32'h7F16C6F4;	13'h02B6: data <= 32'h7F1EE11C;	13'h02B7: data <= 32'h7F26D6B9;	13'h02B8: data <= 32'h7F2EA7C8;	13'h02B9: data <= 32'h7F365448;	13'h02BA: data <= 32'h7F3DDC36;	13'h02BB: data <= 32'h7F453F8F;	13'h02BC: data <= 32'h7F4C7E52;	13'h02BD: data <= 32'h7F53987D;	13'h02BE: data <= 32'h7F5A8E0E;	13'h02BF: data <= 32'h7F615F02;	13'h02C0: data <= 32'h7F680B58;	13'h02C1: data <= 32'h7F6E930E;	13'h02C2: data <= 32'h7F74F622;	13'h02C3: data <= 32'h7F7B3491;	13'h02C4: data <= 32'h7F814E5B;	13'h02C5: data <= 32'h7F87437E;	13'h02C6: data <= 32'h7F8D13F7;	13'h02C7: data <= 32'h7F92BFC5;	13'h02C8: data <= 32'h7F9846E7;	13'h02C9: data <= 32'h7F9DA95B;	13'h02CA: data <= 32'h7FA2E71F;	13'h02CB: data <= 32'h7FA80032;	13'h02CC: data <= 32'h7FACF493;	13'h02CD: data <= 32'h7FB1C43F;	13'h02CE: data <= 32'h7FB66F36;	13'h02CF: data <= 32'h7FBAF576;	13'h02D0: data <= 32'h7FBF56FE;	13'h02D1: data <= 32'h7FC393CD;	13'h02D2: data <= 32'h7FC7ABE1;	13'h02D3: data <= 32'h7FCB9F39;	13'h02D4: data <= 32'h7FCF6DD5;	13'h02D5: data <= 32'h7FD317B3;	13'h02D6: data <= 32'h7FD69CD1;	13'h02D7: data <= 32'h7FD9FD30;	13'h02D8: data <= 32'h7FDD38CE;	13'h02D9: data <= 32'h7FE04FAA;	13'h02DA: data <= 32'h7FE341C2;	13'h02DB: data <= 32'h7FE60F18;	13'h02DC: data <= 32'h7FE8B7A9;	13'h02DD: data <= 32'h7FEB3B74;	13'h02DE: data <= 32'h7FED9A7A;	13'h02DF: data <= 32'h7FEFD4B9;	13'h02E0: data <= 32'h7FF1EA31;	13'h02E1: data <= 32'h7FF3DAE1;	13'h02E2: data <= 32'h7FF5A6C8;	13'h02E3: data <= 32'h7FF74DE7;	13'h02E4: data <= 32'h7FF8D03C;	13'h02E5: data <= 32'h7FFA2DC7;	13'h02E6: data <= 32'h7FFB6688;	13'h02E7: data <= 32'h7FFC7A7F;	13'h02E8: data <= 32'h7FFD69AA;	13'h02E9: data <= 32'h7FFE340B;	13'h02EA: data <= 32'h7FFED9A0;	13'h02EB: data <= 32'h7FFF5A69;	13'h02EC: data <= 32'h7FFFB667;	13'h02ED: data <= 32'h7FFFED99;	13'h02EE: data <= 32'h7FFFFFFF;	13'h02EF: data <= 32'h7FFFED99;	13'h02F0: data <= 32'h7FFFB667;	13'h02F1: data <= 32'h7FFF5A69;	13'h02F2: data <= 32'h7FFED9A0;	13'h02F3: data <= 32'h7FFE340B;	13'h02F4: data <= 32'h7FFD69AA;	13'h02F5: data <= 32'h7FFC7A7F;	13'h02F6: data <= 32'h7FFB6688;	13'h02F7: data <= 32'h7FFA2DC7;	13'h02F8: data <= 32'h7FF8D03C;	13'h02F9: data <= 32'h7FF74DE7;	13'h02FA: data <= 32'h7FF5A6C8;	13'h02FB: data <= 32'h7FF3DAE1;	13'h02FC: data <= 32'h7FF1EA31;	13'h02FD: data <= 32'h7FEFD4B9;	13'h02FE: data <= 32'h7FED9A7A;	13'h02FF: data <= 32'h7FEB3B74;	13'h0300: data <= 32'h7FE8B7A9;	13'h0301: data <= 32'h7FE60F18;	13'h0302: data <= 32'h7FE341C2;	13'h0303: data <= 32'h7FE04FAA;	13'h0304: data <= 32'h7FDD38CE;	13'h0305: data <= 32'h7FD9FD30;	13'h0306: data <= 32'h7FD69CD1;	13'h0307: data <= 32'h7FD317B3;	13'h0308: data <= 32'h7FCF6DD5;	13'h0309: data <= 32'h7FCB9F39;	13'h030A: data <= 32'h7FC7ABE1;	13'h030B: data <= 32'h7FC393CD;	13'h030C: data <= 32'h7FBF56FE;	13'h030D: data <= 32'h7FBAF576;	13'h030E: data <= 32'h7FB66F36;	13'h030F: data <= 32'h7FB1C43F;	13'h0310: data <= 32'h7FACF493;	13'h0311: data <= 32'h7FA80032;	13'h0312: data <= 32'h7FA2E71F;	13'h0313: data <= 32'h7F9DA95B;	13'h0314: data <= 32'h7F9846E7;	13'h0315: data <= 32'h7F92BFC5;	13'h0316: data <= 32'h7F8D13F7;	13'h0317: data <= 32'h7F87437E;	13'h0318: data <= 32'h7F814E5B;	13'h0319: data <= 32'h7F7B3491;	13'h031A: data <= 32'h7F74F622;	13'h031B: data <= 32'h7F6E930E;	13'h031C: data <= 32'h7F680B58;	13'h031D: data <= 32'h7F615F02;	13'h031E: data <= 32'h7F5A8E0E;	13'h031F: data <= 32'h7F53987D;	13'h0320: data <= 32'h7F4C7E52;	13'h0321: data <= 32'h7F453F8F;	13'h0322: data <= 32'h7F3DDC36;	13'h0323: data <= 32'h7F365448;	13'h0324: data <= 32'h7F2EA7C8;	13'h0325: data <= 32'h7F26D6B9;	13'h0326: data <= 32'h7F1EE11C;	13'h0327: data <= 32'h7F16C6F4;	13'h0328: data <= 32'h7F0E8843;	13'h0329: data <= 32'h7F06250C;	13'h032A: data <= 32'h7EFD9D51;	13'h032B: data <= 32'h7EF4F113;	13'h032C: data <= 32'h7EEC2057;	13'h032D: data <= 32'h7EE32B1E;	13'h032E: data <= 32'h7EDA116B;	13'h032F: data <= 32'h7ED0D341;	13'h0330: data <= 32'h7EC770A2;	13'h0331: data <= 32'h7EBDE991;	13'h0332: data <= 32'h7EB43E11;	13'h0333: data <= 32'h7EAA6E24;	13'h0334: data <= 32'h7EA079CD;	13'h0335: data <= 32'h7E96610F;	13'h0336: data <= 32'h7E8C23EE;	13'h0337: data <= 32'h7E81C26B;	13'h0338: data <= 32'h7E773C8B;	13'h0339: data <= 32'h7E6C924F;	13'h033A: data <= 32'h7E61C3BC;	13'h033B: data <= 32'h7E56D0D3;	13'h033C: data <= 32'h7E4BB999;	13'h033D: data <= 32'h7E407E11;	13'h033E: data <= 32'h7E351E3D;	13'h033F: data <= 32'h7E299A21;	13'h0340: data <= 32'h7E1DF1C1;	13'h0341: data <= 32'h7E12251F;	13'h0342: data <= 32'h7E06343F;	13'h0343: data <= 32'h7DFA1F25;	13'h0344: data <= 32'h7DEDE5D4;	13'h0345: data <= 32'h7DE1884F;	13'h0346: data <= 32'h7DD5069A;	13'h0347: data <= 32'h7DC860B9;	13'h0348: data <= 32'h7DBB96AF;	13'h0349: data <= 32'h7DAEA880;	13'h034A: data <= 32'h7DA19630;	13'h034B: data <= 32'h7D945FC2;	13'h034C: data <= 32'h7D87053A;	13'h034D: data <= 32'h7D79869D;	13'h034E: data <= 32'h7D6BE3ED;	13'h034F: data <= 32'h7D5E1D2F;	13'h0350: data <= 32'h7D503267;	13'h0351: data <= 32'h7D422399;	13'h0352: data <= 32'h7D33F0C8;	13'h0353: data <= 32'h7D2599FA;	13'h0354: data <= 32'h7D171F32;	13'h0355: data <= 32'h7D088073;	13'h0356: data <= 32'h7CF9BDC4;	13'h0357: data <= 32'h7CEAD727;	13'h0358: data <= 32'h7CDBCCA0;	13'h0359: data <= 32'h7CCC9E36;	13'h035A: data <= 32'h7CBD4BEA;	13'h035B: data <= 32'h7CADD5C3;	13'h035C: data <= 32'h7C9E3BC4;	13'h035D: data <= 32'h7C8E7DF3;	13'h035E: data <= 32'h7C7E9C53;	13'h035F: data <= 32'h7C6E96E8;	13'h0360: data <= 32'h7C5E6DB9;	13'h0361: data <= 32'h7C4E20C9;	13'h0362: data <= 32'h7C3DB01C;	13'h0363: data <= 32'h7C2D1BB9;	13'h0364: data <= 32'h7C1C63A3;	13'h0365: data <= 32'h7C0B87DF;	13'h0366: data <= 32'h7BFA8873;	13'h0367: data <= 32'h7BE96562;	13'h0368: data <= 32'h7BD81EB3;	13'h0369: data <= 32'h7BC6B469;	13'h036A: data <= 32'h7BB5268A;	13'h036B: data <= 32'h7BA3751C;	13'h036C: data <= 32'h7B91A022;	13'h036D: data <= 32'h7B7FA7A3;	13'h036E: data <= 32'h7B6D8BA2;	13'h036F: data <= 32'h7B5B4C27;	13'h0370: data <= 32'h7B48E935;	13'h0371: data <= 32'h7B3662D2;	13'h0372: data <= 32'h7B23B904;	13'h0373: data <= 32'h7B10EBD0;	13'h0374: data <= 32'h7AFDFB3A;	13'h0375: data <= 32'h7AEAE74A;	13'h0376: data <= 32'h7AD7B003;	13'h0377: data <= 32'h7AC4556C;	13'h0378: data <= 32'h7AB0D78B;	13'h0379: data <= 32'h7A9D3664;	13'h037A: data <= 32'h7A8971FD;	13'h037B: data <= 32'h7A758A5D;	13'h037C: data <= 32'h7A617F89;	13'h037D: data <= 32'h7A4D5186;	13'h037E: data <= 32'h7A39005A;	13'h037F: data <= 32'h7A248C0C;	13'h0380: data <= 32'h7A0FF4A1;	13'h0381: data <= 32'h79FB3A1F;	13'h0382: data <= 32'h79E65C8C;	13'h0383: data <= 32'h79D15BEE;	13'h0384: data <= 32'h79BC384C;	13'h0385: data <= 32'h79A6F1AA;	13'h0386: data <= 32'h7991880F;	13'h0387: data <= 32'h797BFB82;	13'h0388: data <= 32'h79664C09;	13'h0389: data <= 32'h795079A9;	13'h038A: data <= 32'h793A846A;	13'h038B: data <= 32'h79246C50;	13'h038C: data <= 32'h790E3164;	13'h038D: data <= 32'h78F7D3AB;	13'h038E: data <= 32'h78E1532B;	13'h038F: data <= 32'h78CAAFEC;	13'h0390: data <= 32'h78B3E9F3;	13'h0391: data <= 32'h789D0147;	13'h0392: data <= 32'h7885F5EE;	13'h0393: data <= 32'h786EC7F1;	13'h0394: data <= 32'h78577754;	13'h0395: data <= 32'h7840041E;	13'h0396: data <= 32'h78286E58;	13'h0397: data <= 32'h7810B606;	13'h0398: data <= 32'h77F8DB31;	13'h0399: data <= 32'h77E0DDDE;	13'h039A: data <= 32'h77C8BE15;	13'h039B: data <= 32'h77B07BDD;	13'h039C: data <= 32'h7798173C;	13'h039D: data <= 32'h777F903B;	13'h039E: data <= 32'h7766E6DF;	13'h039F: data <= 32'h774E1B2F;	13'h03A0: data <= 32'h77352D34;	13'h03A1: data <= 32'h771C1CF4;	13'h03A2: data <= 32'h7702EA76;	13'h03A3: data <= 32'h76E995C2;	13'h03A4: data <= 32'h76D01EDF;	13'h03A5: data <= 32'h76B685D4;	13'h03A6: data <= 32'h769CCAA8;	13'h03A7: data <= 32'h7682ED64;	13'h03A8: data <= 32'h7668EE0D;	13'h03A9: data <= 32'h764ECCAD;	13'h03AA: data <= 32'h7634894A;	13'h03AB: data <= 32'h761A23EC;	13'h03AC: data <= 32'h75FF9C9A;	13'h03AD: data <= 32'h75E4F35D;	13'h03AE: data <= 32'h75CA283B;	13'h03AF: data <= 32'h75AF3B3D;	13'h03B0: data <= 32'h75942C6A;	13'h03B1: data <= 32'h7578FBCA;	13'h03B2: data <= 32'h755DA965;	13'h03B3: data <= 32'h75423543;	13'h03B4: data <= 32'h75269F6B;	13'h03B5: data <= 32'h750AE7E5;	13'h03B6: data <= 32'h74EF0EBB;	13'h03B7: data <= 32'h74D313F2;	13'h03B8: data <= 32'h74B6F794;	13'h03B9: data <= 32'h749AB9A9;	13'h03BA: data <= 32'h747E5A39;	13'h03BB: data <= 32'h7461D94B;	13'h03BC: data <= 32'h744536E8;	13'h03BD: data <= 32'h74287319;	13'h03BE: data <= 32'h740B8DE5;	13'h03BF: data <= 32'h73EE8756;	13'h03C0: data <= 32'h73D15F72;	13'h03C1: data <= 32'h73B41643;	13'h03C2: data <= 32'h7396ABD1;	13'h03C3: data <= 32'h73792025;	13'h03C4: data <= 32'h735B7346;	13'h03C5: data <= 32'h733DA53E;	13'h03C6: data <= 32'h731FB615;	13'h03C7: data <= 32'h7301A5D4;	13'h03C8: data <= 32'h72E37483;	13'h03C9: data <= 32'h72C5222B;	13'h03CA: data <= 32'h72A6AED5;	13'h03CB: data <= 32'h72881A89;	13'h03CC: data <= 32'h72696551;	13'h03CD: data <= 32'h724A8F35;	13'h03CE: data <= 32'h722B983D;	13'h03CF: data <= 32'h720C8074;	13'h03D0: data <= 32'h71ED47E1;	13'h03D1: data <= 32'h71CDEE8E;	13'h03D2: data <= 32'h71AE7484;	13'h03D3: data <= 32'h718ED9CB;	13'h03D4: data <= 32'h716F1E6E;	13'h03D5: data <= 32'h714F4274;	13'h03D6: data <= 32'h712F45E8;	13'h03D7: data <= 32'h710F28D2;	13'h03D8: data <= 32'h70EEEB3C;	13'h03D9: data <= 32'h70CE8D2F;	13'h03DA: data <= 32'h70AE0EB4;	13'h03DB: data <= 32'h708D6FD4;	13'h03DC: data <= 32'h706CB09A;	13'h03DD: data <= 32'h704BD10D;	13'h03DE: data <= 32'h702AD139;	13'h03DF: data <= 32'h7009B125;	13'h03E0: data <= 32'h6FE870DD;	13'h03E1: data <= 32'h6FC71069;	13'h03E2: data <= 32'h6FA58FD3;	13'h03E3: data <= 32'h6F83EF24;	13'h03E4: data <= 32'h6F622E67;	13'h03E5: data <= 32'h6F404DA4;	13'h03E6: data <= 32'h6F1E4CE6;	13'h03E7: data <= 32'h6EFC2C37;	13'h03E8: data <= 32'h6ED9EBA0;	13'h03E9: data <= 32'h6EB78B2B;	13'h03EA: data <= 32'h6E950AE2;	13'h03EB: data <= 32'h6E726ACF;	13'h03EC: data <= 32'h6E4FAAFC;	13'h03ED: data <= 32'h6E2CCB73;	13'h03EE: data <= 32'h6E09CC3D;	13'h03EF: data <= 32'h6DE6AD66;	13'h03F0: data <= 32'h6DC36EF7;	13'h03F1: data <= 32'h6DA010F9;	13'h03F2: data <= 32'h6D7C9378;	13'h03F3: data <= 32'h6D58F67E;	13'h03F4: data <= 32'h6D353A15;	13'h03F5: data <= 32'h6D115E46;	13'h03F6: data <= 32'h6CED631D;	13'h03F7: data <= 32'h6CC948A3;	13'h03F8: data <= 32'h6CA50EE4;	13'h03F9: data <= 32'h6C80B5E9;	13'h03FA: data <= 32'h6C5C3DBD;	13'h03FB: data <= 32'h6C37A66B;	13'h03FC: data <= 32'h6C12EFFC;	13'h03FD: data <= 32'h6BEE1A7C;	13'h03FE: data <= 32'h6BC925F5;	13'h03FF: data <= 32'h6BA41272;	13'h0400: data <= 32'h6B7EDFFD;	13'h0401: data <= 32'h6B598EA1;	13'h0402: data <= 32'h6B341E69;	13'h0403: data <= 32'h6B0E8F60;	13'h0404: data <= 32'h6AE8E190;	13'h0405: data <= 32'h6AC31504;	13'h0406: data <= 32'h6A9D29C7;	13'h0407: data <= 32'h6A771FE4;	13'h0408: data <= 32'h6A50F766;	13'h0409: data <= 32'h6A2AB058;	13'h040A: data <= 32'h6A044AC5;	13'h040B: data <= 32'h69DDC6B8;	13'h040C: data <= 32'h69B7243B;	13'h040D: data <= 32'h6990635B;	13'h040E: data <= 32'h69698422;	13'h040F: data <= 32'h6942869B;	13'h0410: data <= 32'h691B6AD2;	13'h0411: data <= 32'h68F430D2;	13'h0412: data <= 32'h68CCD8A5;	13'h0413: data <= 32'h68A56259;	13'h0414: data <= 32'h687DCDF7;	13'h0415: data <= 32'h68561B8B;	13'h0416: data <= 32'h682E4B21;	13'h0417: data <= 32'h68065CC4;	13'h0418: data <= 32'h67DE507F;	13'h0419: data <= 32'h67B6265E;	13'h041A: data <= 32'h678DDE6D;	13'h041B: data <= 32'h676578B7;	13'h041C: data <= 32'h673CF548;	13'h041D: data <= 32'h6714542B;	13'h041E: data <= 32'h66EB956C;	13'h041F: data <= 32'h66C2B917;	13'h0420: data <= 32'h6699BF37;	13'h0421: data <= 32'h6670A7D9;	13'h0422: data <= 32'h66477308;	13'h0423: data <= 32'h661E20D0;	13'h0424: data <= 32'h65F4B13D;	13'h0425: data <= 32'h65CB245A;	13'h0426: data <= 32'h65A17A34;	13'h0427: data <= 32'h6577B2D7;	13'h0428: data <= 32'h654DCE4F;	13'h0429: data <= 32'h6523CCA7;	13'h042A: data <= 32'h64F9ADEC;	13'h042B: data <= 32'h64CF722A;	13'h042C: data <= 32'h64A5196D;	13'h042D: data <= 32'h647AA3C2;	13'h042E: data <= 32'h64501133;	13'h042F: data <= 32'h642561CF;	13'h0430: data <= 32'h63FA95A0;	13'h0431: data <= 32'h63CFACB4;	13'h0432: data <= 32'h63A4A716;	13'h0433: data <= 32'h637984D3;	13'h0434: data <= 32'h634E45F8;	13'h0435: data <= 32'h6322EA90;	13'h0436: data <= 32'h62F772A8;	13'h0437: data <= 32'h62CBDE4E;	13'h0438: data <= 32'h62A02D8C;	13'h0439: data <= 32'h62746071;	13'h043A: data <= 32'h62487707;	13'h043B: data <= 32'h621C715D;	13'h043C: data <= 32'h61F04F7F;	13'h043D: data <= 32'h61C41179;	13'h043E: data <= 32'h6197B758;	13'h043F: data <= 32'h616B4129;	13'h0440: data <= 32'h613EAEF8;	13'h0441: data <= 32'h611200D3;	13'h0442: data <= 32'h60E536C6;	13'h0443: data <= 32'h60B850DF;	13'h0444: data <= 32'h608B4F29;	13'h0445: data <= 32'h605E31B3;	13'h0446: data <= 32'h6030F888;	13'h0447: data <= 32'h6003A3B7;	13'h0448: data <= 32'h5FD6334C;	13'h0449: data <= 32'h5FA8A753;	13'h044A: data <= 32'h5F7AFFDB;	13'h044B: data <= 32'h5F4D3CF0;	13'h044C: data <= 32'h5F1F5EA0;	13'h044D: data <= 32'h5EF164F7;	13'h044E: data <= 32'h5EC35003;	13'h044F: data <= 32'h5E951FD1;	13'h0450: data <= 32'h5E66D46E;	13'h0451: data <= 32'h5E386DE9;	13'h0452: data <= 32'h5E09EC4D;	13'h0453: data <= 32'h5DDB4FA9;	13'h0454: data <= 32'h5DAC9809;	13'h0455: data <= 32'h5D7DC57C;	13'h0456: data <= 32'h5D4ED80E;	13'h0457: data <= 32'h5D1FCFCE;	13'h0458: data <= 32'h5CF0ACC8;	13'h0459: data <= 32'h5CC16F0A;	13'h045A: data <= 32'h5C9216A3;	13'h045B: data <= 32'h5C62A39E;	13'h045C: data <= 32'h5C33160B;	13'h045D: data <= 32'h5C036DF7;	13'h045E: data <= 32'h5BD3AB6F;	13'h045F: data <= 32'h5BA3CE81;	13'h0460: data <= 32'h5B73D73B;	13'h0461: data <= 32'h5B43C5AB;	13'h0462: data <= 32'h5B1399DF;	13'h0463: data <= 32'h5AE353E3;	13'h0464: data <= 32'h5AB2F3C7;	13'h0465: data <= 32'h5A827999;	13'h0466: data <= 32'h5A51E565;	13'h0467: data <= 32'h5A21373B;	13'h0468: data <= 32'h59F06F27;	13'h0469: data <= 32'h59BF8D39;	13'h046A: data <= 32'h598E917E;	13'h046B: data <= 32'h595D7C04;	13'h046C: data <= 32'h592C4CD9;	13'h046D: data <= 32'h58FB040C;	13'h046E: data <= 32'h58C9A1AA;	13'h046F: data <= 32'h589825C3;	13'h0470: data <= 32'h58669063;	13'h0471: data <= 32'h5834E19A;	13'h0472: data <= 32'h58031975;	13'h0473: data <= 32'h57D13804;	13'h0474: data <= 32'h579F3D53;	13'h0475: data <= 32'h576D2972;	13'h0476: data <= 32'h573AFC6F;	13'h0477: data <= 32'h5708B659;	13'h0478: data <= 32'h56D6573E;	13'h0479: data <= 32'h56A3DF2B;	13'h047A: data <= 32'h56714E31;	13'h047B: data <= 32'h563EA45D;	13'h047C: data <= 32'h560BE1BF;	13'h047D: data <= 32'h55D90663;	13'h047E: data <= 32'h55A6125A;	13'h047F: data <= 32'h557305B2;	13'h0480: data <= 32'h553FE07A;	13'h0481: data <= 32'h550CA2BF;	13'h0482: data <= 32'h54D94C92;	13'h0483: data <= 32'h54A5DE00;	13'h0484: data <= 32'h54725719;	13'h0485: data <= 32'h543EB7EB;	13'h0486: data <= 32'h540B0085;	13'h0487: data <= 32'h53D730F6;	13'h0488: data <= 32'h53A3494D;	13'h0489: data <= 32'h536F4999;	13'h048A: data <= 32'h533B31E9;	13'h048B: data <= 32'h5307024B;	13'h048C: data <= 32'h52D2BAD0;	13'h048D: data <= 32'h529E5B85;	13'h048E: data <= 32'h5269E47A;	13'h048F: data <= 32'h523555BD;	13'h0490: data <= 32'h5200AF5F;	13'h0491: data <= 32'h51CBF16E;	13'h0492: data <= 32'h51971BFA;	13'h0493: data <= 32'h51622F11;	13'h0494: data <= 32'h512D2AC2;	13'h0495: data <= 32'h50F80F1E;	13'h0496: data <= 32'h50C2DC33;	13'h0497: data <= 32'h508D9210;	13'h0498: data <= 32'h505830C5;	13'h0499: data <= 32'h5022B862;	13'h049A: data <= 32'h4FED28F5;	13'h049B: data <= 32'h4FB7828E;	13'h049C: data <= 32'h4F81C53C;	13'h049D: data <= 32'h4F4BF10F;	13'h049E: data <= 32'h4F160617;	13'h049F: data <= 32'h4EE00462;	13'h04A0: data <= 32'h4EA9EC01;	13'h04A1: data <= 32'h4E73BD02;	13'h04A2: data <= 32'h4E3D7776;	13'h04A3: data <= 32'h4E071B6D;	13'h04A4: data <= 32'h4DD0A8F4;	13'h04A5: data <= 32'h4D9A201D;	13'h04A6: data <= 32'h4D6380F8;	13'h04A7: data <= 32'h4D2CCB93;	13'h04A8: data <= 32'h4CF5FFFE;	13'h04A9: data <= 32'h4CBF1E4A;	13'h04AA: data <= 32'h4C882685;	13'h04AB: data <= 32'h4C5118C0;	13'h04AC: data <= 32'h4C19F50B;	13'h04AD: data <= 32'h4BE2BB76;	13'h04AE: data <= 32'h4BAB6C10;	13'h04AF: data <= 32'h4B7406E9;	13'h04B0: data <= 32'h4B3C8C11;	13'h04B1: data <= 32'h4B04FB98;	13'h04B2: data <= 32'h4ACD558E;	13'h04B3: data <= 32'h4A959A04;	13'h04B4: data <= 32'h4A5DC908;	13'h04B5: data <= 32'h4A25E2AC;	13'h04B6: data <= 32'h49EDE6FF;	13'h04B7: data <= 32'h49B5D611;	13'h04B8: data <= 32'h497DAFF3;	13'h04B9: data <= 32'h494574B4;	13'h04BA: data <= 32'h490D2465;	13'h04BB: data <= 32'h48D4BF16;	13'h04BC: data <= 32'h489C44D7;	13'h04BD: data <= 32'h4863B5B9;	13'h04BE: data <= 32'h482B11CB;	13'h04BF: data <= 32'h47F2591E;	13'h04C0: data <= 32'h47B98BC2;	13'h04C1: data <= 32'h4780A9C8;	13'h04C2: data <= 32'h4747B33F;	13'h04C3: data <= 32'h470EA839;	13'h04C4: data <= 32'h46D588C6;	13'h04C5: data <= 32'h469C54F6;	13'h04C6: data <= 32'h46630CD9;	13'h04C7: data <= 32'h4629B080;	13'h04C8: data <= 32'h45F03FFC;	13'h04C9: data <= 32'h45B6BB5D;	13'h04CA: data <= 32'h457D22B3;	13'h04CB: data <= 32'h4543760F;	13'h04CC: data <= 32'h4509B583;	13'h04CD: data <= 32'h44CFE11D;	13'h04CE: data <= 32'h4495F8EF;	13'h04CF: data <= 32'h445BFD0A;	13'h04D0: data <= 32'h4421ED7E;	13'h04D1: data <= 32'h43E7CA5C;	13'h04D2: data <= 32'h43AD93B5;	13'h04D3: data <= 32'h43734999;	13'h04D4: data <= 32'h4338EC19;	13'h04D5: data <= 32'h42FE7B46;	13'h04D6: data <= 32'h42C3F731;	13'h04D7: data <= 32'h42895FEA;	13'h04D8: data <= 32'h424EB583;	13'h04D9: data <= 32'h4213F80C;	13'h04DA: data <= 32'h41D92796;	13'h04DB: data <= 32'h419E4432;	13'h04DC: data <= 32'h41634DF1;	13'h04DD: data <= 32'h412844E3;	13'h04DE: data <= 32'h40ED291B;	13'h04DF: data <= 32'h40B1FAA9;	13'h04E0: data <= 32'h4076B99D;	13'h04E1: data <= 32'h403B660A;	13'h04E2: data <= 32'h3FFFFFFF;	13'h04E3: data <= 32'h3FC4878E;	13'h04E4: data <= 32'h3F88FCC9;	13'h04E5: data <= 32'h3F4D5FC0;	13'h04E6: data <= 32'h3F11B084;	13'h04E7: data <= 32'h3ED5EF27;	13'h04E8: data <= 32'h3E9A1BB9;	13'h04E9: data <= 32'h3E5E364C;	13'h04EA: data <= 32'h3E223EF2;	13'h04EB: data <= 32'h3DE635BB;	13'h04EC: data <= 32'h3DAA1AB9;	13'h04ED: data <= 32'h3D6DEDFC;	13'h04EE: data <= 32'h3D31AF97;	13'h04EF: data <= 32'h3CF55F9A;	13'h04F0: data <= 32'h3CB8FE17;	13'h04F1: data <= 32'h3C7C8B1F;	13'h04F2: data <= 32'h3C4006C4;	13'h04F3: data <= 32'h3C037117;	13'h04F4: data <= 32'h3BC6CA2A;	13'h04F5: data <= 32'h3B8A120D;	13'h04F6: data <= 32'h3B4D48D3;	13'h04F7: data <= 32'h3B106E8C;	13'h04F8: data <= 32'h3AD3834B;	13'h04F9: data <= 32'h3A968720;	13'h04FA: data <= 32'h3A597A1E;	13'h04FB: data <= 32'h3A1C5C56;	13'h04FC: data <= 32'h39DF2DD9;	13'h04FD: data <= 32'h39A1EEB9;	13'h04FE: data <= 32'h39649F08;	13'h04FF: data <= 32'h39273ED7;	13'h0500: data <= 32'h38E9CE38;	13'h0501: data <= 32'h38AC4D3C;	13'h0502: data <= 32'h386EBBF6;	13'h0503: data <= 32'h38311A77;	13'h0504: data <= 32'h37F368D0;	13'h0505: data <= 32'h37B5A714;	13'h0506: data <= 32'h3777D554;	13'h0507: data <= 32'h3739F3A2;	13'h0508: data <= 32'h36FC0210;	13'h0509: data <= 32'h36BE00AF;	13'h050A: data <= 32'h367FEF91;	13'h050B: data <= 32'h3641CEC9;	13'h050C: data <= 32'h36039E68;	13'h050D: data <= 32'h35C55E80;	13'h050E: data <= 32'h35870F22;	13'h050F: data <= 32'h3548B061;	13'h0510: data <= 32'h350A424F;	13'h0511: data <= 32'h34CBC4FE;	13'h0512: data <= 32'h348D387F;	13'h0513: data <= 32'h344E9CE5;	13'h0514: data <= 32'h340FF241;	13'h0515: data <= 32'h33D138A6;	13'h0516: data <= 32'h33927025;	13'h0517: data <= 32'h335398D2;	13'h0518: data <= 32'h3314B2BC;	13'h0519: data <= 32'h32D5BDF8;	13'h051A: data <= 32'h3296BA97;	13'h051B: data <= 32'h3257A8AA;	13'h051C: data <= 32'h32188845;	13'h051D: data <= 32'h31D95979;	13'h051E: data <= 32'h319A1C58;	13'h051F: data <= 32'h315AD0F5;	13'h0520: data <= 32'h311B7762;	13'h0521: data <= 32'h30DC0FB1;	13'h0522: data <= 32'h309C99F5;	13'h0523: data <= 32'h305D163E;	13'h0524: data <= 32'h301D84A1;	13'h0525: data <= 32'h2FDDE52E;	13'h0526: data <= 32'h2F9E37F9;	13'h0527: data <= 32'h2F5E7D14;	13'h0528: data <= 32'h2F1EB490;	13'h0529: data <= 32'h2EDEDE81;	13'h052A: data <= 32'h2E9EFAF9;	13'h052B: data <= 32'h2E5F0A09;	13'h052C: data <= 32'h2E1F0BC5;	13'h052D: data <= 32'h2DDF003F;	13'h052E: data <= 32'h2D9EE789;	13'h052F: data <= 32'h2D5EC1B5;	13'h0530: data <= 32'h2D1E8ED7;	13'h0531: data <= 32'h2CDE4F00;	13'h0532: data <= 32'h2C9E0243;	13'h0533: data <= 32'h2C5DA8B3;	13'h0534: data <= 32'h2C1D4261;	13'h0535: data <= 32'h2BDCCF61;	13'h0536: data <= 32'h2B9C4FC5;	13'h0537: data <= 32'h2B5BC3A0;	13'h0538: data <= 32'h2B1B2B04;	13'h0539: data <= 32'h2ADA8603;	13'h053A: data <= 32'h2A99D4B1;	13'h053B: data <= 32'h2A59171F;	13'h053C: data <= 32'h2A184D61;	13'h053D: data <= 32'h29D7778A;	13'h053E: data <= 32'h299695AA;	13'h053F: data <= 32'h2955A7D7;	13'h0540: data <= 32'h2914AE21;	13'h0541: data <= 32'h28D3A89C;	13'h0542: data <= 32'h2892975B;	13'h0543: data <= 32'h28517A6F;	13'h0544: data <= 32'h281051ED;	13'h0545: data <= 32'h27CF1DE6;	13'h0546: data <= 32'h278DDE6E;	13'h0547: data <= 32'h274C9396;	13'h0548: data <= 32'h270B3D72;	13'h0549: data <= 32'h26C9DC16;	13'h054A: data <= 32'h26886F92;	13'h054B: data <= 32'h2646F7FB;	13'h054C: data <= 32'h26057562;	13'h054D: data <= 32'h25C3E7DC;	13'h054E: data <= 32'h25824F7A;	13'h054F: data <= 32'h2540AC50;	13'h0550: data <= 32'h24FEFE71;	13'h0551: data <= 32'h24BD45EF;	13'h0552: data <= 32'h247B82DD;	13'h0553: data <= 32'h2439B54E;	13'h0554: data <= 32'h23F7DD55;	13'h0555: data <= 32'h23B5FB05;	13'h0556: data <= 32'h23740E72;	13'h0557: data <= 32'h233217AD;	13'h0558: data <= 32'h22F016C9;	13'h0559: data <= 32'h22AE0BDB;	13'h055A: data <= 32'h226BF6F5;	13'h055B: data <= 32'h2229D829;	13'h055C: data <= 32'h21E7AF8B;	13'h055D: data <= 32'h21A57D2E;	13'h055E: data <= 32'h21634125;	13'h055F: data <= 32'h2120FB82;	13'h0560: data <= 32'h20DEAC5A;	13'h0561: data <= 32'h209C53BF;	13'h0562: data <= 32'h2059F1C3;	13'h0563: data <= 32'h2017867B;	13'h0564: data <= 32'h1FD511F9;	13'h0565: data <= 32'h1F929451;	13'h0566: data <= 32'h1F500D95;	13'h0567: data <= 32'h1F0D7DD8;	13'h0568: data <= 32'h1ECAE52F;	13'h0569: data <= 32'h1E8843AB;	13'h056A: data <= 32'h1E459960;	13'h056B: data <= 32'h1E02E662;	13'h056C: data <= 32'h1DC02AC2;	13'h056D: data <= 32'h1D7D6696;	13'h056E: data <= 32'h1D3A99EF;	13'h056F: data <= 32'h1CF7C4E1;	13'h0570: data <= 32'h1CB4E77F;	13'h0571: data <= 32'h1C7201DD;	13'h0572: data <= 32'h1C2F140D;	13'h0573: data <= 32'h1BEC1E23;	13'h0574: data <= 32'h1BA92032;	13'h0575: data <= 32'h1B661A4E;	13'h0576: data <= 32'h1B230C89;	13'h0577: data <= 32'h1ADFF6F7;	13'h0578: data <= 32'h1A9CD9AC;	13'h0579: data <= 32'h1A59B4B9;	13'h057A: data <= 32'h1A168834;	13'h057B: data <= 32'h19D3542F;	13'h057C: data <= 32'h199018BD;	13'h057D: data <= 32'h194CD5F2;	13'h057E: data <= 32'h19098BE1;	13'h057F: data <= 32'h18C63A9D;	13'h0580: data <= 32'h1882E23A;	13'h0581: data <= 32'h183F82CC;	13'h0582: data <= 32'h17FC1C64;	13'h0583: data <= 32'h17B8AF18;	13'h0584: data <= 32'h17753AFA;	13'h0585: data <= 32'h1731C01E;	13'h0586: data <= 32'h16EE3E96;	13'h0587: data <= 32'h16AAB677;	13'h0588: data <= 32'h166727D4;	13'h0589: data <= 32'h162392C1;	13'h058A: data <= 32'h15DFF750;	13'h058B: data <= 32'h159C5595;	13'h058C: data <= 32'h1558ADA4;	13'h058D: data <= 32'h1514FF90;	13'h058E: data <= 32'h14D14B6C;	13'h058F: data <= 32'h148D914D;	13'h0590: data <= 32'h1449D144;	13'h0591: data <= 32'h14060B67;	13'h0592: data <= 32'h13C23FC8;	13'h0593: data <= 32'h137E6E7B;	13'h0594: data <= 32'h133A9793;	13'h0595: data <= 32'h12F6BB25;	13'h0596: data <= 32'h12B2D942;	13'h0597: data <= 32'h126EF200;	13'h0598: data <= 32'h122B0571;	13'h0599: data <= 32'h11E713A9;	13'h059A: data <= 32'h11A31CBB;	13'h059B: data <= 32'h115F20BC;	13'h059C: data <= 32'h111B1FBE;	13'h059D: data <= 32'h10D719D5;	13'h059E: data <= 32'h10930F15;	13'h059F: data <= 32'h104EFF91;	13'h05A0: data <= 32'h100AEB5D;	13'h05A1: data <= 32'h0FC6D28C;	13'h05A2: data <= 32'h0F82B532;	13'h05A3: data <= 32'h0F3E9363;	13'h05A4: data <= 32'h0EFA6D32;	13'h05A5: data <= 32'h0EB642B3;	13'h05A6: data <= 32'h0E7213F8;	13'h05A7: data <= 32'h0E2DE117;	13'h05A8: data <= 32'h0DE9AA23;	13'h05A9: data <= 32'h0DA56F2E;	13'h05AA: data <= 32'h0D61304D;	13'h05AB: data <= 32'h0D1CED93;	13'h05AC: data <= 32'h0CD8A715;	13'h05AD: data <= 32'h0C945CE5;	13'h05AE: data <= 32'h0C500F17;	13'h05AF: data <= 32'h0C0BBDBF;	13'h05B0: data <= 32'h0BC768F1;	13'h05B1: data <= 32'h0B8310C0;	13'h05B2: data <= 32'h0B3EB53F;	13'h05B3: data <= 32'h0AFA5684;	13'h05B4: data <= 32'h0AB5F4A0;	13'h05B5: data <= 32'h0A718FA8;	13'h05B6: data <= 32'h0A2D27AF;	13'h05B7: data <= 32'h09E8BCC9;	13'h05B8: data <= 32'h09A44F0B;	13'h05B9: data <= 32'h095FDE86;	13'h05BA: data <= 32'h091B6B50;	13'h05BB: data <= 32'h08D6F57B;	13'h05BC: data <= 32'h08927D1C;	13'h05BD: data <= 32'h084E0246;	13'h05BE: data <= 32'h0809850D;	13'h05BF: data <= 32'h07C50585;	13'h05C0: data <= 32'h078083C0;	13'h05C1: data <= 32'h073BFFD4;	13'h05C2: data <= 32'h06F779D3;	13'h05C3: data <= 32'h06B2F1D2;	13'h05C4: data <= 32'h066E67E3;	13'h05C5: data <= 32'h0629DC1B;	13'h05C6: data <= 32'h05E54E8E;	13'h05C7: data <= 32'h05A0BF4F;	13'h05C8: data <= 32'h055C2E71;	13'h05C9: data <= 32'h05179C09;	13'h05CA: data <= 32'h04D3082A;	13'h05CB: data <= 32'h048E72E9;	13'h05CC: data <= 32'h0449DC58;	13'h05CD: data <= 32'h0405448B;	13'h05CE: data <= 32'h03C0AB96;	13'h05CF: data <= 32'h037C118E;	13'h05D0: data <= 32'h03377685;	13'h05D1: data <= 32'h02F2DA8F;	13'h05D2: data <= 32'h02AE3DC0;	13'h05D3: data <= 32'h0269A02C;	13'h05D4: data <= 32'h022501E6;	13'h05D5: data <= 32'h01E06302;	13'h05D6: data <= 32'h019BC395;	13'h05D7: data <= 32'h015723B1;	13'h05D8: data <= 32'h0112836A;	13'h05D9: data <= 32'h00CDE2D4;	13'h05DA: data <= 32'h00894204;	13'h05DB: data <= 32'h0044A10B;	13'h05DC: data <= 32'h00000000;	13'h05DD: data <= 32'hFFBB5EF5;	13'h05DE: data <= 32'hFF76BDFC;	13'h05DF: data <= 32'hFF321D2C;	13'h05E0: data <= 32'hFEED7C96;	13'h05E1: data <= 32'hFEA8DC4F;	13'h05E2: data <= 32'hFE643C6B;	13'h05E3: data <= 32'hFE1F9CFE;	13'h05E4: data <= 32'hFDDAFE1A;	13'h05E5: data <= 32'hFD965FD4;	13'h05E6: data <= 32'hFD51C240;	13'h05E7: data <= 32'hFD0D2571;	13'h05E8: data <= 32'hFCC8897B;	13'h05E9: data <= 32'hFC83EE72;	13'h05EA: data <= 32'hFC3F546A;	13'h05EB: data <= 32'hFBFABB75;	13'h05EC: data <= 32'hFBB623A8;	13'h05ED: data <= 32'hFB718D17;	13'h05EE: data <= 32'hFB2CF7D6;	13'h05EF: data <= 32'hFAE863F7;	13'h05F0: data <= 32'hFAA3D18F;	13'h05F1: data <= 32'hFA5F40B1;	13'h05F2: data <= 32'hFA1AB172;	13'h05F3: data <= 32'hF9D623E5;	13'h05F4: data <= 32'hF991981D;	13'h05F5: data <= 32'hF94D0E2E;	13'h05F6: data <= 32'hF908862D;	13'h05F7: data <= 32'hF8C4002C;	13'h05F8: data <= 32'hF87F7C40;	13'h05F9: data <= 32'hF83AFA7B;	13'h05FA: data <= 32'hF7F67AF3;	13'h05FB: data <= 32'hF7B1FDBA;	13'h05FC: data <= 32'hF76D82E4;	13'h05FD: data <= 32'hF7290A85;	13'h05FE: data <= 32'hF6E494B0;	13'h05FF: data <= 32'hF6A0217A;	13'h0600: data <= 32'hF65BB0F5;	13'h0601: data <= 32'hF6174337;	13'h0602: data <= 32'hF5D2D851;	13'h0603: data <= 32'hF58E7058;	13'h0604: data <= 32'hF54A0B60;	13'h0605: data <= 32'hF505A97C;	13'h0606: data <= 32'hF4C14AC1;	13'h0607: data <= 32'hF47CEF40;	13'h0608: data <= 32'hF438970F;	13'h0609: data <= 32'hF3F44241;	13'h060A: data <= 32'hF3AFF0E9;	13'h060B: data <= 32'hF36BA31B;	13'h060C: data <= 32'hF32758EB;	13'h060D: data <= 32'hF2E3126D;	13'h060E: data <= 32'hF29ECFB3;	13'h060F: data <= 32'hF25A90D2;	13'h0610: data <= 32'hF21655DD;	13'h0611: data <= 32'hF1D21EE9;	13'h0612: data <= 32'hF18DEC08;	13'h0613: data <= 32'hF149BD4D;	13'h0614: data <= 32'hF10592CE;	13'h0615: data <= 32'hF0C16C9D;	13'h0616: data <= 32'hF07D4ACE;	13'h0617: data <= 32'hF0392D74;	13'h0618: data <= 32'hEFF514A3;	13'h0619: data <= 32'hEFB1006F;	13'h061A: data <= 32'hEF6CF0EB;	13'h061B: data <= 32'hEF28E62B;	13'h061C: data <= 32'hEEE4E042;	13'h061D: data <= 32'hEEA0DF44;	13'h061E: data <= 32'hEE5CE345;	13'h061F: data <= 32'hEE18EC57;	13'h0620: data <= 32'hEDD4FA8F;	13'h0621: data <= 32'hED910E00;	13'h0622: data <= 32'hED4D26BE;	13'h0623: data <= 32'hED0944DB;	13'h0624: data <= 32'hECC5686D;	13'h0625: data <= 32'hEC819185;	13'h0626: data <= 32'hEC3DC038;	13'h0627: data <= 32'hEBF9F499;	13'h0628: data <= 32'hEBB62EBC;	13'h0629: data <= 32'hEB726EB3;	13'h062A: data <= 32'hEB2EB494;	13'h062B: data <= 32'hEAEB0070;	13'h062C: data <= 32'hEAA7525C;	13'h062D: data <= 32'hEA63AA6B;	13'h062E: data <= 32'hEA2008B0;	13'h062F: data <= 32'hE9DC6D3F;	13'h0630: data <= 32'hE998D82C;	13'h0631: data <= 32'hE9554989;	13'h0632: data <= 32'hE911C16A;	13'h0633: data <= 32'hE8CE3FE2;	13'h0634: data <= 32'hE88AC506;	13'h0635: data <= 32'hE84750E8;	13'h0636: data <= 32'hE803E39C;	13'h0637: data <= 32'hE7C07D34;	13'h0638: data <= 32'hE77D1DC6;	13'h0639: data <= 32'hE739C563;	13'h063A: data <= 32'hE6F6741F;	13'h063B: data <= 32'hE6B32A0E;	13'h063C: data <= 32'hE66FE743;	13'h063D: data <= 32'hE62CABD1;	13'h063E: data <= 32'hE5E977CC;	13'h063F: data <= 32'hE5A64B47;	13'h0640: data <= 32'hE5632654;	13'h0641: data <= 32'hE5200909;	13'h0642: data <= 32'hE4DCF377;	13'h0643: data <= 32'hE499E5B2;	13'h0644: data <= 32'hE456DFCE;	13'h0645: data <= 32'hE413E1DD;	13'h0646: data <= 32'hE3D0EBF3;	13'h0647: data <= 32'hE38DFE23;	13'h0648: data <= 32'hE34B1881;	13'h0649: data <= 32'hE3083B1F;	13'h064A: data <= 32'hE2C56611;	13'h064B: data <= 32'hE282996A;	13'h064C: data <= 32'hE23FD53E;	13'h064D: data <= 32'hE1FD199E;	13'h064E: data <= 32'hE1BA66A0;	13'h064F: data <= 32'hE177BC55;	13'h0650: data <= 32'hE1351AD1;	13'h0651: data <= 32'hE0F28228;	13'h0652: data <= 32'hE0AFF26B;	13'h0653: data <= 32'hE06D6BAF;	13'h0654: data <= 32'hE02AEE07;	13'h0655: data <= 32'hDFE87985;	13'h0656: data <= 32'hDFA60E3D;	13'h0657: data <= 32'hDF63AC41;	13'h0658: data <= 32'hDF2153A6;	13'h0659: data <= 32'hDEDF047E;	13'h065A: data <= 32'hDE9CBEDB;	13'h065B: data <= 32'hDE5A82D2;	13'h065C: data <= 32'hDE185075;	13'h065D: data <= 32'hDDD627D7;	13'h065E: data <= 32'hDD94090B;	13'h065F: data <= 32'hDD51F425;	13'h0660: data <= 32'hDD0FE937;	13'h0661: data <= 32'hDCCDE853;	13'h0662: data <= 32'hDC8BF18E;	13'h0663: data <= 32'hDC4A04FB;	13'h0664: data <= 32'hDC0822AB;	13'h0665: data <= 32'hDBC64AB2;	13'h0666: data <= 32'hDB847D23;	13'h0667: data <= 32'hDB42BA11;	13'h0668: data <= 32'hDB01018F;	13'h0669: data <= 32'hDABF53B0;	13'h066A: data <= 32'hDA7DB086;	13'h066B: data <= 32'hDA3C1824;	13'h066C: data <= 32'hD9FA8A9E;	13'h066D: data <= 32'hD9B90805;	13'h066E: data <= 32'hD977906E;	13'h066F: data <= 32'hD93623EA;	13'h0670: data <= 32'hD8F4C28E;	13'h0671: data <= 32'hD8B36C6A;	13'h0672: data <= 32'hD8722192;	13'h0673: data <= 32'hD830E21A;	13'h0674: data <= 32'hD7EFAE13;	13'h0675: data <= 32'hD7AE8591;	13'h0676: data <= 32'hD76D68A5;	13'h0677: data <= 32'hD72C5764;	13'h0678: data <= 32'hD6EB51DF;	13'h0679: data <= 32'hD6AA5829;	13'h067A: data <= 32'hD6696A56;	13'h067B: data <= 32'hD6288876;	13'h067C: data <= 32'hD5E7B29F;	13'h067D: data <= 32'hD5A6E8E1;	13'h067E: data <= 32'hD5662B4F;	13'h067F: data <= 32'hD52579FD;	13'h0680: data <= 32'hD4E4D4FC;	13'h0681: data <= 32'hD4A43C60;	13'h0682: data <= 32'hD463B03B;	13'h0683: data <= 32'hD423309F;	13'h0684: data <= 32'hD3E2BD9F;	13'h0685: data <= 32'hD3A2574D;	13'h0686: data <= 32'hD361FDBD;	13'h0687: data <= 32'hD321B100;	13'h0688: data <= 32'hD2E17129;	13'h0689: data <= 32'hD2A13E4B;	13'h068A: data <= 32'hD2611877;	13'h068B: data <= 32'hD220FFC1;	13'h068C: data <= 32'hD1E0F43B;	13'h068D: data <= 32'hD1A0F5F7;	13'h068E: data <= 32'hD1610507;	13'h068F: data <= 32'hD121217F;	13'h0690: data <= 32'hD0E14B70;	13'h0691: data <= 32'hD0A182EC;	13'h0692: data <= 32'hD061C807;	13'h0693: data <= 32'hD0221AD2;	13'h0694: data <= 32'hCFE27B5F;	13'h0695: data <= 32'hCFA2E9C2;	13'h0696: data <= 32'hCF63660B;	13'h0697: data <= 32'hCF23F04F;	13'h0698: data <= 32'hCEE4889E;	13'h0699: data <= 32'hCEA52F0B;	13'h069A: data <= 32'hCE65E3A8;	13'h069B: data <= 32'hCE26A687;	13'h069C: data <= 32'hCDE777BB;	13'h069D: data <= 32'hCDA85756;	13'h069E: data <= 32'hCD694569;	13'h069F: data <= 32'hCD2A4208;	13'h06A0: data <= 32'hCCEB4D44;	13'h06A1: data <= 32'hCCAC672E;	13'h06A2: data <= 32'hCC6D8FDB;	13'h06A3: data <= 32'hCC2EC75A;	13'h06A4: data <= 32'hCBF00DBF;	13'h06A5: data <= 32'hCBB1631B;	13'h06A6: data <= 32'hCB72C781;	13'h06A7: data <= 32'hCB343B02;	13'h06A8: data <= 32'hCAF5BDB1;	13'h06A9: data <= 32'hCAB74F9F;	13'h06AA: data <= 32'hCA78F0DE;	13'h06AB: data <= 32'hCA3AA180;	13'h06AC: data <= 32'hC9FC6198;	13'h06AD: data <= 32'hC9BE3137;	13'h06AE: data <= 32'hC980106F;	13'h06AF: data <= 32'hC941FF51;	13'h06B0: data <= 32'hC903FDF0;	13'h06B1: data <= 32'hC8C60C5E;	13'h06B2: data <= 32'hC8882AAC;	13'h06B3: data <= 32'hC84A58EC;	13'h06B4: data <= 32'hC80C9730;	13'h06B5: data <= 32'hC7CEE589;	13'h06B6: data <= 32'hC791440A;	13'h06B7: data <= 32'hC753B2C4;	13'h06B8: data <= 32'hC71631C8;	13'h06B9: data <= 32'hC6D8C129;	13'h06BA: data <= 32'hC69B60F8;	13'h06BB: data <= 32'hC65E1147;	13'h06BC: data <= 32'hC620D227;	13'h06BD: data <= 32'hC5E3A3AA;	13'h06BE: data <= 32'hC5A685E2;	13'h06BF: data <= 32'hC56978E0;	13'h06C0: data <= 32'hC52C7CB5;	13'h06C1: data <= 32'hC4EF9174;	13'h06C2: data <= 32'hC4B2B72D;	13'h06C3: data <= 32'hC475EDF3;	13'h06C4: data <= 32'hC43935D6;	13'h06C5: data <= 32'hC3FC8EE9;	13'h06C6: data <= 32'hC3BFF93C;	13'h06C7: data <= 32'hC38374E1;	13'h06C8: data <= 32'hC34701E9;	13'h06C9: data <= 32'hC30AA066;	13'h06CA: data <= 32'hC2CE5069;	13'h06CB: data <= 32'hC2921204;	13'h06CC: data <= 32'hC255E547;	13'h06CD: data <= 32'hC219CA45;	13'h06CE: data <= 32'hC1DDC10E;	13'h06CF: data <= 32'hC1A1C9B4;	13'h06D0: data <= 32'hC165E447;	13'h06D1: data <= 32'hC12A10D9;	13'h06D2: data <= 32'hC0EE4F7C;	13'h06D3: data <= 32'hC0B2A040;	13'h06D4: data <= 32'hC0770337;	13'h06D5: data <= 32'hC03B7872;	13'h06D6: data <= 32'hC0000001;	13'h06D7: data <= 32'hBFC499F6;	13'h06D8: data <= 32'hBF894663;	13'h06D9: data <= 32'hBF4E0557;	13'h06DA: data <= 32'hBF12D6E5;	13'h06DB: data <= 32'hBED7BB1D;	13'h06DC: data <= 32'hBE9CB20F;	13'h06DD: data <= 32'hBE61BBCE;	13'h06DE: data <= 32'hBE26D86A;	13'h06DF: data <= 32'hBDEC07F4;	13'h06E0: data <= 32'hBDB14A7D;	13'h06E1: data <= 32'hBD76A016;	13'h06E2: data <= 32'hBD3C08CF;	13'h06E3: data <= 32'hBD0184BA;	13'h06E4: data <= 32'hBCC713E7;	13'h06E5: data <= 32'hBC8CB667;	13'h06E6: data <= 32'hBC526C4B;	13'h06E7: data <= 32'hBC1835A4;	13'h06E8: data <= 32'hBBDE1282;	13'h06E9: data <= 32'hBBA402F6;	13'h06EA: data <= 32'hBB6A0711;	13'h06EB: data <= 32'hBB301EE3;	13'h06EC: data <= 32'hBAF64A7D;	13'h06ED: data <= 32'hBABC89F1;	13'h06EE: data <= 32'hBA82DD4D;	13'h06EF: data <= 32'hBA4944A3;	13'h06F0: data <= 32'hBA0FC004;	13'h06F1: data <= 32'hB9D64F80;	13'h06F2: data <= 32'hB99CF327;	13'h06F3: data <= 32'hB963AB0A;	13'h06F4: data <= 32'hB92A773A;	13'h06F5: data <= 32'hB8F157C7;	13'h06F6: data <= 32'hB8B84CC1;	13'h06F7: data <= 32'hB87F5638;	13'h06F8: data <= 32'hB846743E;	13'h06F9: data <= 32'hB80DA6E2;	13'h06FA: data <= 32'hB7D4EE35;	13'h06FB: data <= 32'hB79C4A47;	13'h06FC: data <= 32'hB763BB29;	13'h06FD: data <= 32'hB72B40EA;	13'h06FE: data <= 32'hB6F2DB9B;	13'h06FF: data <= 32'hB6BA8B4C;	13'h0700: data <= 32'hB682500D;	13'h0701: data <= 32'hB64A29EF;	13'h0702: data <= 32'hB6121901;	13'h0703: data <= 32'hB5DA1D54;	13'h0704: data <= 32'hB5A236F8;	13'h0705: data <= 32'hB56A65FC;	13'h0706: data <= 32'hB532AA72;	13'h0707: data <= 32'hB4FB0468;	13'h0708: data <= 32'hB4C373EF;	13'h0709: data <= 32'hB48BF917;	13'h070A: data <= 32'hB45493F0;	13'h070B: data <= 32'hB41D448A;	13'h070C: data <= 32'hB3E60AF5;	13'h070D: data <= 32'hB3AEE740;	13'h070E: data <= 32'hB377D97B;	13'h070F: data <= 32'hB340E1B6;	13'h0710: data <= 32'hB30A0002;	13'h0711: data <= 32'hB2D3346D;	13'h0712: data <= 32'hB29C7F08;	13'h0713: data <= 32'hB265DFE3;	13'h0714: data <= 32'hB22F570C;	13'h0715: data <= 32'hB1F8E493;	13'h0716: data <= 32'hB1C2888A;	13'h0717: data <= 32'hB18C42FE;	13'h0718: data <= 32'hB15613FF;	13'h0719: data <= 32'hB11FFB9E;	13'h071A: data <= 32'hB0E9F9E9;	13'h071B: data <= 32'hB0B40EF1;	13'h071C: data <= 32'hB07E3AC4;	13'h071D: data <= 32'hB0487D72;	13'h071E: data <= 32'hB012D70B;	13'h071F: data <= 32'hAFDD479E;	13'h0720: data <= 32'hAFA7CF3B;	13'h0721: data <= 32'hAF726DF0;	13'h0722: data <= 32'hAF3D23CD;	13'h0723: data <= 32'hAF07F0E2;	13'h0724: data <= 32'hAED2D53E;	13'h0725: data <= 32'hAE9DD0EF;	13'h0726: data <= 32'hAE68E406;	13'h0727: data <= 32'hAE340E92;	13'h0728: data <= 32'hADFF50A1;	13'h0729: data <= 32'hADCAAA43;	13'h072A: data <= 32'hAD961B86;	13'h072B: data <= 32'hAD61A47B;	13'h072C: data <= 32'hAD2D4530;	13'h072D: data <= 32'hACF8FDB5;	13'h072E: data <= 32'hACC4CE17;	13'h072F: data <= 32'hAC90B667;	13'h0730: data <= 32'hAC5CB6B3;	13'h0731: data <= 32'hAC28CF0A;	13'h0732: data <= 32'hABF4FF7B;	13'h0733: data <= 32'hABC14815;	13'h0734: data <= 32'hAB8DA8E7;	13'h0735: data <= 32'hAB5A2200;	13'h0736: data <= 32'hAB26B36E;	13'h0737: data <= 32'hAAF35D41;	13'h0738: data <= 32'hAAC01F86;	13'h0739: data <= 32'hAA8CFA4E;	13'h073A: data <= 32'hAA59EDA6;	13'h073B: data <= 32'hAA26F99D;	13'h073C: data <= 32'hA9F41E41;	13'h073D: data <= 32'hA9C15BA3;	13'h073E: data <= 32'hA98EB1CF;	13'h073F: data <= 32'hA95C20D5;	13'h0740: data <= 32'hA929A8C2;	13'h0741: data <= 32'hA8F749A7;	13'h0742: data <= 32'hA8C50391;	13'h0743: data <= 32'hA892D68E;	13'h0744: data <= 32'hA860C2AD;	13'h0745: data <= 32'hA82EC7FC;	13'h0746: data <= 32'hA7FCE68B;	13'h0747: data <= 32'hA7CB1E66;	13'h0748: data <= 32'hA7996F9D;	13'h0749: data <= 32'hA767DA3D;	13'h074A: data <= 32'hA7365E56;	13'h074B: data <= 32'hA704FBF4;	13'h074C: data <= 32'hA6D3B327;	13'h074D: data <= 32'hA6A283FC;	13'h074E: data <= 32'hA6716E82;	13'h074F: data <= 32'hA64072C7;	13'h0750: data <= 32'hA60F90D9;	13'h0751: data <= 32'hA5DEC8C5;	13'h0752: data <= 32'hA5AE1A9B;	13'h0753: data <= 32'hA57D8667;	13'h0754: data <= 32'hA54D0C39;	13'h0755: data <= 32'hA51CAC1D;	13'h0756: data <= 32'hA4EC6621;	13'h0757: data <= 32'hA4BC3A55;	13'h0758: data <= 32'hA48C28C5;	13'h0759: data <= 32'hA45C317F;	13'h075A: data <= 32'hA42C5491;	13'h075B: data <= 32'hA3FC9209;	13'h075C: data <= 32'hA3CCE9F5;	13'h075D: data <= 32'hA39D5C62;	13'h075E: data <= 32'hA36DE95D;	13'h075F: data <= 32'hA33E90F6;	13'h0760: data <= 32'hA30F5338;	13'h0761: data <= 32'hA2E03032;	13'h0762: data <= 32'hA2B127F2;	13'h0763: data <= 32'hA2823A84;	13'h0764: data <= 32'hA25367F7;	13'h0765: data <= 32'hA224B057;	13'h0766: data <= 32'hA1F613B3;	13'h0767: data <= 32'hA1C79217;	13'h0768: data <= 32'hA1992B92;	13'h0769: data <= 32'hA16AE02F;	13'h076A: data <= 32'hA13CAFFD;	13'h076B: data <= 32'hA10E9B09;	13'h076C: data <= 32'hA0E0A160;	13'h076D: data <= 32'hA0B2C310;	13'h076E: data <= 32'hA0850025;	13'h076F: data <= 32'hA05758AD;	13'h0770: data <= 32'hA029CCB4;	13'h0771: data <= 32'h9FFC5C49;	13'h0772: data <= 32'h9FCF0778;	13'h0773: data <= 32'h9FA1CE4D;	13'h0774: data <= 32'h9F74B0D7;	13'h0775: data <= 32'h9F47AF21;	13'h0776: data <= 32'h9F1AC93A;	13'h0777: data <= 32'h9EEDFF2D;	13'h0778: data <= 32'h9EC15108;	13'h0779: data <= 32'h9E94BED7;	13'h077A: data <= 32'h9E6848A8;	13'h077B: data <= 32'h9E3BEE87;	13'h077C: data <= 32'h9E0FB081;	13'h077D: data <= 32'h9DE38EA3;	13'h077E: data <= 32'h9DB788F9;	13'h077F: data <= 32'h9D8B9F8F;	13'h0780: data <= 32'h9D5FD274;	13'h0781: data <= 32'h9D3421B2;	13'h0782: data <= 32'h9D088D58;	13'h0783: data <= 32'h9CDD1570;	13'h0784: data <= 32'h9CB1BA08;	13'h0785: data <= 32'h9C867B2D;	13'h0786: data <= 32'h9C5B58EA;	13'h0787: data <= 32'h9C30534C;	13'h0788: data <= 32'h9C056A60;	13'h0789: data <= 32'h9BDA9E31;	13'h078A: data <= 32'h9BAFEECD;	13'h078B: data <= 32'h9B855C3E;	13'h078C: data <= 32'h9B5AE693;	13'h078D: data <= 32'h9B308DD6;	13'h078E: data <= 32'h9B065214;	13'h078F: data <= 32'h9ADC3359;	13'h0790: data <= 32'h9AB231B1;	13'h0791: data <= 32'h9A884D29;	13'h0792: data <= 32'h9A5E85CC;	13'h0793: data <= 32'h9A34DBA6;	13'h0794: data <= 32'h9A0B4EC3;	13'h0795: data <= 32'h99E1DF30;	13'h0796: data <= 32'h99B88CF8;	13'h0797: data <= 32'h998F5827;	13'h0798: data <= 32'h996640C9;	13'h0799: data <= 32'h993D46E9;	13'h079A: data <= 32'h99146A94;	13'h079B: data <= 32'h98EBABD5;	13'h079C: data <= 32'h98C30AB8;	13'h079D: data <= 32'h989A8749;	13'h079E: data <= 32'h98722193;	13'h079F: data <= 32'h9849D9A2;	13'h07A0: data <= 32'h9821AF81;	13'h07A1: data <= 32'h97F9A33C;	13'h07A2: data <= 32'h97D1B4DF;	13'h07A3: data <= 32'h97A9E475;	13'h07A4: data <= 32'h97823209;	13'h07A5: data <= 32'h975A9DA7;	13'h07A6: data <= 32'h9733275B;	13'h07A7: data <= 32'h970BCF2E;	13'h07A8: data <= 32'h96E4952E;	13'h07A9: data <= 32'h96BD7965;	13'h07AA: data <= 32'h96967BDE;	13'h07AB: data <= 32'h966F9CA5;	13'h07AC: data <= 32'h9648DBC5;	13'h07AD: data <= 32'h96223948;	13'h07AE: data <= 32'h95FBB53B;	13'h07AF: data <= 32'h95D54FA8;	13'h07B0: data <= 32'h95AF089A;	13'h07B1: data <= 32'h9588E01C;	13'h07B2: data <= 32'h9562D639;	13'h07B3: data <= 32'h953CEAFC;	13'h07B4: data <= 32'h95171E70;	13'h07B5: data <= 32'h94F170A0;	13'h07B6: data <= 32'h94CBE197;	13'h07B7: data <= 32'h94A6715F;	13'h07B8: data <= 32'h94812003;	13'h07B9: data <= 32'h945BED8E;	13'h07BA: data <= 32'h9436DA0B;	13'h07BB: data <= 32'h9411E584;	13'h07BC: data <= 32'h93ED1004;	13'h07BD: data <= 32'h93C85995;	13'h07BE: data <= 32'h93A3C243;	13'h07BF: data <= 32'h937F4A17;	13'h07C0: data <= 32'h935AF11C;	13'h07C1: data <= 32'h9336B75D;	13'h07C2: data <= 32'h93129CE3;	13'h07C3: data <= 32'h92EEA1BA;	13'h07C4: data <= 32'h92CAC5EB;	13'h07C5: data <= 32'h92A70982;	13'h07C6: data <= 32'h92836C88;	13'h07C7: data <= 32'h925FEF07;	13'h07C8: data <= 32'h923C9109;	13'h07C9: data <= 32'h9219529A;	13'h07CA: data <= 32'h91F633C3;	13'h07CB: data <= 32'h91D3348D;	13'h07CC: data <= 32'h91B05504;	13'h07CD: data <= 32'h918D9531;	13'h07CE: data <= 32'h916AF51E;	13'h07CF: data <= 32'h914874D5;	13'h07D0: data <= 32'h91261460;	13'h07D1: data <= 32'h9103D3C9;	13'h07D2: data <= 32'h90E1B31A;	13'h07D3: data <= 32'h90BFB25C;	13'h07D4: data <= 32'h909DD199;	13'h07D5: data <= 32'h907C10DC;	13'h07D6: data <= 32'h905A702D;	13'h07D7: data <= 32'h9038EF97;	13'h07D8: data <= 32'h90178F23;	13'h07D9: data <= 32'h8FF64EDB;	13'h07DA: data <= 32'h8FD52EC7;	13'h07DB: data <= 32'h8FB42EF3;	13'h07DC: data <= 32'h8F934F66;	13'h07DD: data <= 32'h8F72902C;	13'h07DE: data <= 32'h8F51F14C;	13'h07DF: data <= 32'h8F3172D1;	13'h07E0: data <= 32'h8F1114C4;	13'h07E1: data <= 32'h8EF0D72E;	13'h07E2: data <= 32'h8ED0BA18;	13'h07E3: data <= 32'h8EB0BD8C;	13'h07E4: data <= 32'h8E90E192;	13'h07E5: data <= 32'h8E712635;	13'h07E6: data <= 32'h8E518B7C;	13'h07E7: data <= 32'h8E321172;	13'h07E8: data <= 32'h8E12B81F;	13'h07E9: data <= 32'h8DF37F8C;	13'h07EA: data <= 32'h8DD467C3;	13'h07EB: data <= 32'h8DB570CB;	13'h07EC: data <= 32'h8D969AAF;	13'h07ED: data <= 32'h8D77E577;	13'h07EE: data <= 32'h8D59512B;	13'h07EF: data <= 32'h8D3ADDD5;	13'h07F0: data <= 32'h8D1C8B7D;	13'h07F1: data <= 32'h8CFE5A2C;	13'h07F2: data <= 32'h8CE049EB;	13'h07F3: data <= 32'h8CC25AC2;	13'h07F4: data <= 32'h8CA48CBA;	13'h07F5: data <= 32'h8C86DFDB;	13'h07F6: data <= 32'h8C69542F;	13'h07F7: data <= 32'h8C4BE9BD;	13'h07F8: data <= 32'h8C2EA08E;	13'h07F9: data <= 32'h8C1178AA;	13'h07FA: data <= 32'h8BF4721B;	13'h07FB: data <= 32'h8BD78CE7;	13'h07FC: data <= 32'h8BBAC918;	13'h07FD: data <= 32'h8B9E26B5;	13'h07FE: data <= 32'h8B81A5C7;	13'h07FF: data <= 32'h8B654657;	13'h0800: data <= 32'h8B49086C;	13'h0801: data <= 32'h8B2CEC0E;	13'h0802: data <= 32'h8B10F145;	13'h0803: data <= 32'h8AF5181B;	13'h0804: data <= 32'h8AD96095;	13'h0805: data <= 32'h8ABDCABD;	13'h0806: data <= 32'h8AA2569B;	13'h0807: data <= 32'h8A870436;	13'h0808: data <= 32'h8A6BD396;	13'h0809: data <= 32'h8A50C4C3;	13'h080A: data <= 32'h8A35D7C5;	13'h080B: data <= 32'h8A1B0CA3;	13'h080C: data <= 32'h8A006366;	13'h080D: data <= 32'h89E5DC14;	13'h080E: data <= 32'h89CB76B6;	13'h080F: data <= 32'h89B13353;	13'h0810: data <= 32'h899711F3;	13'h0811: data <= 32'h897D129C;	13'h0812: data <= 32'h89633558;	13'h0813: data <= 32'h89497A2C;	13'h0814: data <= 32'h892FE121;	13'h0815: data <= 32'h89166A3E;	13'h0816: data <= 32'h88FD158A;	13'h0817: data <= 32'h88E3E30C;	13'h0818: data <= 32'h88CAD2CC;	13'h0819: data <= 32'h88B1E4D1;	13'h081A: data <= 32'h88991921;	13'h081B: data <= 32'h88806FC5;	13'h081C: data <= 32'h8867E8C4;	13'h081D: data <= 32'h884F8423;	13'h081E: data <= 32'h883741EB;	13'h081F: data <= 32'h881F2222;	13'h0820: data <= 32'h880724CF;	13'h0821: data <= 32'h87EF49FA;	13'h0822: data <= 32'h87D791A8;	13'h0823: data <= 32'h87BFFBE2;	13'h0824: data <= 32'h87A888AC;	13'h0825: data <= 32'h8791380F;	13'h0826: data <= 32'h877A0A12;	13'h0827: data <= 32'h8762FEB9;	13'h0828: data <= 32'h874C160D;	13'h0829: data <= 32'h87355014;	13'h082A: data <= 32'h871EACD5;	13'h082B: data <= 32'h87082C55;	13'h082C: data <= 32'h86F1CE9C;	13'h082D: data <= 32'h86DB93B0;	13'h082E: data <= 32'h86C57B96;	13'h082F: data <= 32'h86AF8657;	13'h0830: data <= 32'h8699B3F7;	13'h0831: data <= 32'h8684047E;	13'h0832: data <= 32'h866E77F1;	13'h0833: data <= 32'h86590E56;	13'h0834: data <= 32'h8643C7B4;	13'h0835: data <= 32'h862EA412;	13'h0836: data <= 32'h8619A374;	13'h0837: data <= 32'h8604C5E1;	13'h0838: data <= 32'h85F00B5F;	13'h0839: data <= 32'h85DB73F4;	13'h083A: data <= 32'h85C6FFA6;	13'h083B: data <= 32'h85B2AE7A;	13'h083C: data <= 32'h859E8077;	13'h083D: data <= 32'h858A75A3;	13'h083E: data <= 32'h85768E03;	13'h083F: data <= 32'h8562C99C;	13'h0840: data <= 32'h854F2875;	13'h0841: data <= 32'h853BAA94;	13'h0842: data <= 32'h85284FFD;	13'h0843: data <= 32'h851518B6;	13'h0844: data <= 32'h850204C6;	13'h0845: data <= 32'h84EF1430;	13'h0846: data <= 32'h84DC46FC;	13'h0847: data <= 32'h84C99D2E;	13'h0848: data <= 32'h84B716CB;	13'h0849: data <= 32'h84A4B3D9;	13'h084A: data <= 32'h8492745E;	13'h084B: data <= 32'h8480585D;	13'h084C: data <= 32'h846E5FDE;	13'h084D: data <= 32'h845C8AE4;	13'h084E: data <= 32'h844AD976;	13'h084F: data <= 32'h84394B97;	13'h0850: data <= 32'h8427E14D;	13'h0851: data <= 32'h84169A9E;	13'h0852: data <= 32'h8405778D;	13'h0853: data <= 32'h83F47821;	13'h0854: data <= 32'h83E39C5D;	13'h0855: data <= 32'h83D2E447;	13'h0856: data <= 32'h83C24FE4;	13'h0857: data <= 32'h83B1DF37;	13'h0858: data <= 32'h83A19247;	13'h0859: data <= 32'h83916918;	13'h085A: data <= 32'h838163AD;	13'h085B: data <= 32'h8371820D;	13'h085C: data <= 32'h8361C43C;	13'h085D: data <= 32'h83522A3D;	13'h085E: data <= 32'h8342B416;	13'h085F: data <= 32'h833361CA;	13'h0860: data <= 32'h83243360;	13'h0861: data <= 32'h831528D9;	13'h0862: data <= 32'h8306423C;	13'h0863: data <= 32'h82F77F8D;	13'h0864: data <= 32'h82E8E0CE;	13'h0865: data <= 32'h82DA6606;	13'h0866: data <= 32'h82CC0F38;	13'h0867: data <= 32'h82BDDC67;	13'h0868: data <= 32'h82AFCD99;	13'h0869: data <= 32'h82A1E2D1;	13'h086A: data <= 32'h82941C13;	13'h086B: data <= 32'h82867963;	13'h086C: data <= 32'h8278FAC6;	13'h086D: data <= 32'h826BA03E;	13'h086E: data <= 32'h825E69D0;	13'h086F: data <= 32'h82515780;	13'h0870: data <= 32'h82446951;	13'h0871: data <= 32'h82379F47;	13'h0872: data <= 32'h822AF966;	13'h0873: data <= 32'h821E77B1;	13'h0874: data <= 32'h82121A2C;	13'h0875: data <= 32'h8205E0DB;	13'h0876: data <= 32'h81F9CBC1;	13'h0877: data <= 32'h81EDDAE1;	13'h0878: data <= 32'h81E20E3F;	13'h0879: data <= 32'h81D665DF;	13'h087A: data <= 32'h81CAE1C3;	13'h087B: data <= 32'h81BF81EF;	13'h087C: data <= 32'h81B44667;	13'h087D: data <= 32'h81A92F2D;	13'h087E: data <= 32'h819E3C44;	13'h087F: data <= 32'h81936DB1;	13'h0880: data <= 32'h8188C375;	13'h0881: data <= 32'h817E3D95;	13'h0882: data <= 32'h8173DC12;	13'h0883: data <= 32'h81699EF1;	13'h0884: data <= 32'h815F8633;	13'h0885: data <= 32'h815591DC;	13'h0886: data <= 32'h814BC1EF;	13'h0887: data <= 32'h8142166F;	13'h0888: data <= 32'h81388F5E;	13'h0889: data <= 32'h812F2CBF;	13'h088A: data <= 32'h8125EE95;	13'h088B: data <= 32'h811CD4E2;	13'h088C: data <= 32'h8113DFA9;	13'h088D: data <= 32'h810B0EED;	13'h088E: data <= 32'h810262AF;	13'h088F: data <= 32'h80F9DAF4;	13'h0890: data <= 32'h80F177BD;	13'h0891: data <= 32'h80E9390C;	13'h0892: data <= 32'h80E11EE4;	13'h0893: data <= 32'h80D92947;	13'h0894: data <= 32'h80D15838;	13'h0895: data <= 32'h80C9ABB8;	13'h0896: data <= 32'h80C223CA;	13'h0897: data <= 32'h80BAC071;	13'h0898: data <= 32'h80B381AE;	13'h0899: data <= 32'h80AC6783;	13'h089A: data <= 32'h80A571F2;	13'h089B: data <= 32'h809EA0FE;	13'h089C: data <= 32'h8097F4A8;	13'h089D: data <= 32'h80916CF2;	13'h089E: data <= 32'h808B09DE;	13'h089F: data <= 32'h8084CB6F;	13'h08A0: data <= 32'h807EB1A5;	13'h08A1: data <= 32'h8078BC82;	13'h08A2: data <= 32'h8072EC09;	13'h08A3: data <= 32'h806D403B;	13'h08A4: data <= 32'h8067B919;	13'h08A5: data <= 32'h806256A5;	13'h08A6: data <= 32'h805D18E1;	13'h08A7: data <= 32'h8057FFCE;	13'h08A8: data <= 32'h80530B6D;	13'h08A9: data <= 32'h804E3BC1;	13'h08AA: data <= 32'h804990CA;	13'h08AB: data <= 32'h80450A8A;	13'h08AC: data <= 32'h8040A902;	13'h08AD: data <= 32'h803C6C33;	13'h08AE: data <= 32'h8038541F;	13'h08AF: data <= 32'h803460C7;	13'h08B0: data <= 32'h8030922B;	13'h08B1: data <= 32'h802CE84D;	13'h08B2: data <= 32'h8029632F;	13'h08B3: data <= 32'h802602D0;	13'h08B4: data <= 32'h8022C732;	13'h08B5: data <= 32'h801FB056;	13'h08B6: data <= 32'h801CBE3E;	13'h08B7: data <= 32'h8019F0E8;	13'h08B8: data <= 32'h80174857;	13'h08B9: data <= 32'h8014C48C;	13'h08BA: data <= 32'h80126586;	13'h08BB: data <= 32'h80102B47;	13'h08BC: data <= 32'h800E15CF;	13'h08BD: data <= 32'h800C251F;	13'h08BE: data <= 32'h800A5938;	13'h08BF: data <= 32'h8008B219;	13'h08C0: data <= 32'h80072FC4;	13'h08C1: data <= 32'h8005D239;	13'h08C2: data <= 32'h80049978;	13'h08C3: data <= 32'h80038581;	13'h08C4: data <= 32'h80029656;	13'h08C5: data <= 32'h8001CBF5;	13'h08C6: data <= 32'h80012660;	13'h08C7: data <= 32'h8000A597;	13'h08C8: data <= 32'h80004999;	13'h08C9: data <= 32'h80001267;	13'h08CA: data <= 32'h80000001;	13'h08CB: data <= 32'h80001267;	13'h08CC: data <= 32'h80004999;	13'h08CD: data <= 32'h8000A597;	13'h08CE: data <= 32'h80012660;	13'h08CF: data <= 32'h8001CBF5;	13'h08D0: data <= 32'h80029656;	13'h08D1: data <= 32'h80038581;	13'h08D2: data <= 32'h80049978;	13'h08D3: data <= 32'h8005D239;	13'h08D4: data <= 32'h80072FC4;	13'h08D5: data <= 32'h8008B219;	13'h08D6: data <= 32'h800A5938;	13'h08D7: data <= 32'h800C251F;	13'h08D8: data <= 32'h800E15CF;	13'h08D9: data <= 32'h80102B47;	13'h08DA: data <= 32'h80126586;	13'h08DB: data <= 32'h8014C48C;	13'h08DC: data <= 32'h80174857;	13'h08DD: data <= 32'h8019F0E8;	13'h08DE: data <= 32'h801CBE3E;	13'h08DF: data <= 32'h801FB056;	13'h08E0: data <= 32'h8022C732;	13'h08E1: data <= 32'h802602D0;	13'h08E2: data <= 32'h8029632F;	13'h08E3: data <= 32'h802CE84D;	13'h08E4: data <= 32'h8030922B;	13'h08E5: data <= 32'h803460C7;	13'h08E6: data <= 32'h8038541F;	13'h08E7: data <= 32'h803C6C33;	13'h08E8: data <= 32'h8040A902;	13'h08E9: data <= 32'h80450A8A;	13'h08EA: data <= 32'h804990CA;	13'h08EB: data <= 32'h804E3BC1;	13'h08EC: data <= 32'h80530B6D;	13'h08ED: data <= 32'h8057FFCE;	13'h08EE: data <= 32'h805D18E1;	13'h08EF: data <= 32'h806256A5;	13'h08F0: data <= 32'h8067B919;	13'h08F1: data <= 32'h806D403B;	13'h08F2: data <= 32'h8072EC09;	13'h08F3: data <= 32'h8078BC82;	13'h08F4: data <= 32'h807EB1A5;	13'h08F5: data <= 32'h8084CB6F;	13'h08F6: data <= 32'h808B09DE;	13'h08F7: data <= 32'h80916CF2;	13'h08F8: data <= 32'h8097F4A8;	13'h08F9: data <= 32'h809EA0FE;	13'h08FA: data <= 32'h80A571F2;	13'h08FB: data <= 32'h80AC6783;	13'h08FC: data <= 32'h80B381AE;	13'h08FD: data <= 32'h80BAC071;	13'h08FE: data <= 32'h80C223CA;	13'h08FF: data <= 32'h80C9ABB8;	13'h0900: data <= 32'h80D15838;	13'h0901: data <= 32'h80D92947;	13'h0902: data <= 32'h80E11EE4;	13'h0903: data <= 32'h80E9390C;	13'h0904: data <= 32'h80F177BD;	13'h0905: data <= 32'h80F9DAF4;	13'h0906: data <= 32'h810262AF;	13'h0907: data <= 32'h810B0EED;	13'h0908: data <= 32'h8113DFA9;	13'h0909: data <= 32'h811CD4E2;	13'h090A: data <= 32'h8125EE95;	13'h090B: data <= 32'h812F2CBF;	13'h090C: data <= 32'h81388F5E;	13'h090D: data <= 32'h8142166F;	13'h090E: data <= 32'h814BC1EF;	13'h090F: data <= 32'h815591DC;	13'h0910: data <= 32'h815F8633;	13'h0911: data <= 32'h81699EF1;	13'h0912: data <= 32'h8173DC12;	13'h0913: data <= 32'h817E3D95;	13'h0914: data <= 32'h8188C375;	13'h0915: data <= 32'h81936DB1;	13'h0916: data <= 32'h819E3C44;	13'h0917: data <= 32'h81A92F2D;	13'h0918: data <= 32'h81B44667;	13'h0919: data <= 32'h81BF81EF;	13'h091A: data <= 32'h81CAE1C3;	13'h091B: data <= 32'h81D665DF;	13'h091C: data <= 32'h81E20E3F;	13'h091D: data <= 32'h81EDDAE1;	13'h091E: data <= 32'h81F9CBC1;	13'h091F: data <= 32'h8205E0DB;	13'h0920: data <= 32'h82121A2C;	13'h0921: data <= 32'h821E77B1;	13'h0922: data <= 32'h822AF966;	13'h0923: data <= 32'h82379F47;	13'h0924: data <= 32'h82446951;	13'h0925: data <= 32'h82515780;	13'h0926: data <= 32'h825E69D0;	13'h0927: data <= 32'h826BA03E;	13'h0928: data <= 32'h8278FAC6;	13'h0929: data <= 32'h82867963;	13'h092A: data <= 32'h82941C13;	13'h092B: data <= 32'h82A1E2D1;	13'h092C: data <= 32'h82AFCD99;	13'h092D: data <= 32'h82BDDC67;	13'h092E: data <= 32'h82CC0F38;	13'h092F: data <= 32'h82DA6606;	13'h0930: data <= 32'h82E8E0CE;	13'h0931: data <= 32'h82F77F8D;	13'h0932: data <= 32'h8306423C;	13'h0933: data <= 32'h831528D9;	13'h0934: data <= 32'h83243360;	13'h0935: data <= 32'h833361CA;	13'h0936: data <= 32'h8342B416;	13'h0937: data <= 32'h83522A3D;	13'h0938: data <= 32'h8361C43C;	13'h0939: data <= 32'h8371820D;	13'h093A: data <= 32'h838163AD;	13'h093B: data <= 32'h83916918;	13'h093C: data <= 32'h83A19247;	13'h093D: data <= 32'h83B1DF37;	13'h093E: data <= 32'h83C24FE4;	13'h093F: data <= 32'h83D2E447;	13'h0940: data <= 32'h83E39C5D;	13'h0941: data <= 32'h83F47821;	13'h0942: data <= 32'h8405778D;	13'h0943: data <= 32'h84169A9E;	13'h0944: data <= 32'h8427E14D;	13'h0945: data <= 32'h84394B97;	13'h0946: data <= 32'h844AD976;	13'h0947: data <= 32'h845C8AE4;	13'h0948: data <= 32'h846E5FDE;	13'h0949: data <= 32'h8480585D;	13'h094A: data <= 32'h8492745E;	13'h094B: data <= 32'h84A4B3D9;	13'h094C: data <= 32'h84B716CB;	13'h094D: data <= 32'h84C99D2E;	13'h094E: data <= 32'h84DC46FC;	13'h094F: data <= 32'h84EF1430;	13'h0950: data <= 32'h850204C6;	13'h0951: data <= 32'h851518B6;	13'h0952: data <= 32'h85284FFD;	13'h0953: data <= 32'h853BAA94;	13'h0954: data <= 32'h854F2875;	13'h0955: data <= 32'h8562C99C;	13'h0956: data <= 32'h85768E03;	13'h0957: data <= 32'h858A75A3;	13'h0958: data <= 32'h859E8077;	13'h0959: data <= 32'h85B2AE7A;	13'h095A: data <= 32'h85C6FFA6;	13'h095B: data <= 32'h85DB73F4;	13'h095C: data <= 32'h85F00B5F;	13'h095D: data <= 32'h8604C5E1;	13'h095E: data <= 32'h8619A374;	13'h095F: data <= 32'h862EA412;	13'h0960: data <= 32'h8643C7B4;	13'h0961: data <= 32'h86590E56;	13'h0962: data <= 32'h866E77F1;	13'h0963: data <= 32'h8684047E;	13'h0964: data <= 32'h8699B3F7;	13'h0965: data <= 32'h86AF8657;	13'h0966: data <= 32'h86C57B96;	13'h0967: data <= 32'h86DB93B0;	13'h0968: data <= 32'h86F1CE9C;	13'h0969: data <= 32'h87082C55;	13'h096A: data <= 32'h871EACD5;	13'h096B: data <= 32'h87355014;	13'h096C: data <= 32'h874C160D;	13'h096D: data <= 32'h8762FEB9;	13'h096E: data <= 32'h877A0A12;	13'h096F: data <= 32'h8791380F;	13'h0970: data <= 32'h87A888AC;	13'h0971: data <= 32'h87BFFBE2;	13'h0972: data <= 32'h87D791A8;	13'h0973: data <= 32'h87EF49FA;	13'h0974: data <= 32'h880724CF;	13'h0975: data <= 32'h881F2222;	13'h0976: data <= 32'h883741EB;	13'h0977: data <= 32'h884F8423;	13'h0978: data <= 32'h8867E8C4;	13'h0979: data <= 32'h88806FC5;	13'h097A: data <= 32'h88991921;	13'h097B: data <= 32'h88B1E4D1;	13'h097C: data <= 32'h88CAD2CC;	13'h097D: data <= 32'h88E3E30C;	13'h097E: data <= 32'h88FD158A;	13'h097F: data <= 32'h89166A3E;	13'h0980: data <= 32'h892FE121;	13'h0981: data <= 32'h89497A2C;	13'h0982: data <= 32'h89633558;	13'h0983: data <= 32'h897D129C;	13'h0984: data <= 32'h899711F3;	13'h0985: data <= 32'h89B13353;	13'h0986: data <= 32'h89CB76B6;	13'h0987: data <= 32'h89E5DC14;	13'h0988: data <= 32'h8A006366;	13'h0989: data <= 32'h8A1B0CA3;	13'h098A: data <= 32'h8A35D7C5;	13'h098B: data <= 32'h8A50C4C3;	13'h098C: data <= 32'h8A6BD396;	13'h098D: data <= 32'h8A870436;	13'h098E: data <= 32'h8AA2569B;	13'h098F: data <= 32'h8ABDCABD;	13'h0990: data <= 32'h8AD96095;	13'h0991: data <= 32'h8AF5181B;	13'h0992: data <= 32'h8B10F145;	13'h0993: data <= 32'h8B2CEC0E;	13'h0994: data <= 32'h8B49086C;	13'h0995: data <= 32'h8B654657;	13'h0996: data <= 32'h8B81A5C7;	13'h0997: data <= 32'h8B9E26B5;	13'h0998: data <= 32'h8BBAC918;	13'h0999: data <= 32'h8BD78CE7;	13'h099A: data <= 32'h8BF4721B;	13'h099B: data <= 32'h8C1178AA;	13'h099C: data <= 32'h8C2EA08E;	13'h099D: data <= 32'h8C4BE9BD;	13'h099E: data <= 32'h8C69542F;	13'h099F: data <= 32'h8C86DFDB;	13'h09A0: data <= 32'h8CA48CBA;	13'h09A1: data <= 32'h8CC25AC2;	13'h09A2: data <= 32'h8CE049EB;	13'h09A3: data <= 32'h8CFE5A2C;	13'h09A4: data <= 32'h8D1C8B7D;	13'h09A5: data <= 32'h8D3ADDD5;	13'h09A6: data <= 32'h8D59512B;	13'h09A7: data <= 32'h8D77E577;	13'h09A8: data <= 32'h8D969AAF;	13'h09A9: data <= 32'h8DB570CB;	13'h09AA: data <= 32'h8DD467C3;	13'h09AB: data <= 32'h8DF37F8C;	13'h09AC: data <= 32'h8E12B81F;	13'h09AD: data <= 32'h8E321172;	13'h09AE: data <= 32'h8E518B7C;	13'h09AF: data <= 32'h8E712635;	13'h09B0: data <= 32'h8E90E192;	13'h09B1: data <= 32'h8EB0BD8C;	13'h09B2: data <= 32'h8ED0BA18;	13'h09B3: data <= 32'h8EF0D72E;	13'h09B4: data <= 32'h8F1114C4;	13'h09B5: data <= 32'h8F3172D1;	13'h09B6: data <= 32'h8F51F14C;	13'h09B7: data <= 32'h8F72902C;	13'h09B8: data <= 32'h8F934F66;	13'h09B9: data <= 32'h8FB42EF3;	13'h09BA: data <= 32'h8FD52EC7;	13'h09BB: data <= 32'h8FF64EDB;	13'h09BC: data <= 32'h90178F23;	13'h09BD: data <= 32'h9038EF97;	13'h09BE: data <= 32'h905A702D;	13'h09BF: data <= 32'h907C10DC;	13'h09C0: data <= 32'h909DD199;	13'h09C1: data <= 32'h90BFB25C;	13'h09C2: data <= 32'h90E1B31A;	13'h09C3: data <= 32'h9103D3C9;	13'h09C4: data <= 32'h91261460;	13'h09C5: data <= 32'h914874D5;	13'h09C6: data <= 32'h916AF51E;	13'h09C7: data <= 32'h918D9531;	13'h09C8: data <= 32'h91B05504;	13'h09C9: data <= 32'h91D3348D;	13'h09CA: data <= 32'h91F633C3;	13'h09CB: data <= 32'h9219529A;	13'h09CC: data <= 32'h923C9109;	13'h09CD: data <= 32'h925FEF07;	13'h09CE: data <= 32'h92836C88;	13'h09CF: data <= 32'h92A70982;	13'h09D0: data <= 32'h92CAC5EB;	13'h09D1: data <= 32'h92EEA1BA;	13'h09D2: data <= 32'h93129CE3;	13'h09D3: data <= 32'h9336B75D;	13'h09D4: data <= 32'h935AF11C;	13'h09D5: data <= 32'h937F4A17;	13'h09D6: data <= 32'h93A3C243;	13'h09D7: data <= 32'h93C85995;	13'h09D8: data <= 32'h93ED1004;	13'h09D9: data <= 32'h9411E584;	13'h09DA: data <= 32'h9436DA0B;	13'h09DB: data <= 32'h945BED8E;	13'h09DC: data <= 32'h94812003;	13'h09DD: data <= 32'h94A6715F;	13'h09DE: data <= 32'h94CBE197;	13'h09DF: data <= 32'h94F170A0;	13'h09E0: data <= 32'h95171E70;	13'h09E1: data <= 32'h953CEAFC;	13'h09E2: data <= 32'h9562D639;	13'h09E3: data <= 32'h9588E01C;	13'h09E4: data <= 32'h95AF089A;	13'h09E5: data <= 32'h95D54FA8;	13'h09E6: data <= 32'h95FBB53B;	13'h09E7: data <= 32'h96223948;	13'h09E8: data <= 32'h9648DBC5;	13'h09E9: data <= 32'h966F9CA5;	13'h09EA: data <= 32'h96967BDE;	13'h09EB: data <= 32'h96BD7965;	13'h09EC: data <= 32'h96E4952E;	13'h09ED: data <= 32'h970BCF2E;	13'h09EE: data <= 32'h9733275B;	13'h09EF: data <= 32'h975A9DA7;	13'h09F0: data <= 32'h97823209;	13'h09F1: data <= 32'h97A9E475;	13'h09F2: data <= 32'h97D1B4DF;	13'h09F3: data <= 32'h97F9A33C;	13'h09F4: data <= 32'h9821AF81;	13'h09F5: data <= 32'h9849D9A2;	13'h09F6: data <= 32'h98722193;	13'h09F7: data <= 32'h989A8749;	13'h09F8: data <= 32'h98C30AB8;	13'h09F9: data <= 32'h98EBABD5;	13'h09FA: data <= 32'h99146A94;	13'h09FB: data <= 32'h993D46E9;	13'h09FC: data <= 32'h996640C9;	13'h09FD: data <= 32'h998F5827;	13'h09FE: data <= 32'h99B88CF8;	13'h09FF: data <= 32'h99E1DF30;	13'h0A00: data <= 32'h9A0B4EC3;	13'h0A01: data <= 32'h9A34DBA6;	13'h0A02: data <= 32'h9A5E85CC;	13'h0A03: data <= 32'h9A884D29;	13'h0A04: data <= 32'h9AB231B1;	13'h0A05: data <= 32'h9ADC3359;	13'h0A06: data <= 32'h9B065214;	13'h0A07: data <= 32'h9B308DD6;	13'h0A08: data <= 32'h9B5AE693;	13'h0A09: data <= 32'h9B855C3E;	13'h0A0A: data <= 32'h9BAFEECD;	13'h0A0B: data <= 32'h9BDA9E31;	13'h0A0C: data <= 32'h9C056A60;	13'h0A0D: data <= 32'h9C30534C;	13'h0A0E: data <= 32'h9C5B58EA;	13'h0A0F: data <= 32'h9C867B2D;	13'h0A10: data <= 32'h9CB1BA08;	13'h0A11: data <= 32'h9CDD1570;	13'h0A12: data <= 32'h9D088D58;	13'h0A13: data <= 32'h9D3421B2;	13'h0A14: data <= 32'h9D5FD274;	13'h0A15: data <= 32'h9D8B9F8F;	13'h0A16: data <= 32'h9DB788F9;	13'h0A17: data <= 32'h9DE38EA3;	13'h0A18: data <= 32'h9E0FB081;	13'h0A19: data <= 32'h9E3BEE87;	13'h0A1A: data <= 32'h9E6848A8;	13'h0A1B: data <= 32'h9E94BED7;	13'h0A1C: data <= 32'h9EC15108;	13'h0A1D: data <= 32'h9EEDFF2D;	13'h0A1E: data <= 32'h9F1AC93A;	13'h0A1F: data <= 32'h9F47AF21;	13'h0A20: data <= 32'h9F74B0D7;	13'h0A21: data <= 32'h9FA1CE4D;	13'h0A22: data <= 32'h9FCF0778;	13'h0A23: data <= 32'h9FFC5C49;	13'h0A24: data <= 32'hA029CCB4;	13'h0A25: data <= 32'hA05758AD;	13'h0A26: data <= 32'hA0850025;	13'h0A27: data <= 32'hA0B2C310;	13'h0A28: data <= 32'hA0E0A160;	13'h0A29: data <= 32'hA10E9B09;	13'h0A2A: data <= 32'hA13CAFFD;	13'h0A2B: data <= 32'hA16AE02F;	13'h0A2C: data <= 32'hA1992B92;	13'h0A2D: data <= 32'hA1C79217;	13'h0A2E: data <= 32'hA1F613B3;	13'h0A2F: data <= 32'hA224B057;	13'h0A30: data <= 32'hA25367F7;	13'h0A31: data <= 32'hA2823A84;	13'h0A32: data <= 32'hA2B127F2;	13'h0A33: data <= 32'hA2E03032;	13'h0A34: data <= 32'hA30F5338;	13'h0A35: data <= 32'hA33E90F6;	13'h0A36: data <= 32'hA36DE95D;	13'h0A37: data <= 32'hA39D5C62;	13'h0A38: data <= 32'hA3CCE9F5;	13'h0A39: data <= 32'hA3FC9209;	13'h0A3A: data <= 32'hA42C5491;	13'h0A3B: data <= 32'hA45C317F;	13'h0A3C: data <= 32'hA48C28C5;	13'h0A3D: data <= 32'hA4BC3A55;	13'h0A3E: data <= 32'hA4EC6621;	13'h0A3F: data <= 32'hA51CAC1D;	13'h0A40: data <= 32'hA54D0C39;	13'h0A41: data <= 32'hA57D8667;	13'h0A42: data <= 32'hA5AE1A9B;	13'h0A43: data <= 32'hA5DEC8C5;	13'h0A44: data <= 32'hA60F90D9;	13'h0A45: data <= 32'hA64072C7;	13'h0A46: data <= 32'hA6716E82;	13'h0A47: data <= 32'hA6A283FC;	13'h0A48: data <= 32'hA6D3B327;	13'h0A49: data <= 32'hA704FBF4;	13'h0A4A: data <= 32'hA7365E56;	13'h0A4B: data <= 32'hA767DA3D;	13'h0A4C: data <= 32'hA7996F9D;	13'h0A4D: data <= 32'hA7CB1E66;	13'h0A4E: data <= 32'hA7FCE68B;	13'h0A4F: data <= 32'hA82EC7FC;	13'h0A50: data <= 32'hA860C2AD;	13'h0A51: data <= 32'hA892D68E;	13'h0A52: data <= 32'hA8C50391;	13'h0A53: data <= 32'hA8F749A7;	13'h0A54: data <= 32'hA929A8C2;	13'h0A55: data <= 32'hA95C20D5;	13'h0A56: data <= 32'hA98EB1CF;	13'h0A57: data <= 32'hA9C15BA3;	13'h0A58: data <= 32'hA9F41E41;	13'h0A59: data <= 32'hAA26F99D;	13'h0A5A: data <= 32'hAA59EDA6;	13'h0A5B: data <= 32'hAA8CFA4E;	13'h0A5C: data <= 32'hAAC01F86;	13'h0A5D: data <= 32'hAAF35D41;	13'h0A5E: data <= 32'hAB26B36E;	13'h0A5F: data <= 32'hAB5A2200;	13'h0A60: data <= 32'hAB8DA8E7;	13'h0A61: data <= 32'hABC14815;	13'h0A62: data <= 32'hABF4FF7B;	13'h0A63: data <= 32'hAC28CF0A;	13'h0A64: data <= 32'hAC5CB6B3;	13'h0A65: data <= 32'hAC90B667;	13'h0A66: data <= 32'hACC4CE17;	13'h0A67: data <= 32'hACF8FDB5;	13'h0A68: data <= 32'hAD2D4530;	13'h0A69: data <= 32'hAD61A47B;	13'h0A6A: data <= 32'hAD961B86;	13'h0A6B: data <= 32'hADCAAA43;	13'h0A6C: data <= 32'hADFF50A1;	13'h0A6D: data <= 32'hAE340E92;	13'h0A6E: data <= 32'hAE68E406;	13'h0A6F: data <= 32'hAE9DD0EF;	13'h0A70: data <= 32'hAED2D53E;	13'h0A71: data <= 32'hAF07F0E2;	13'h0A72: data <= 32'hAF3D23CD;	13'h0A73: data <= 32'hAF726DF0;	13'h0A74: data <= 32'hAFA7CF3B;	13'h0A75: data <= 32'hAFDD479E;	13'h0A76: data <= 32'hB012D70B;	13'h0A77: data <= 32'hB0487D72;	13'h0A78: data <= 32'hB07E3AC4;	13'h0A79: data <= 32'hB0B40EF1;	13'h0A7A: data <= 32'hB0E9F9E9;	13'h0A7B: data <= 32'hB11FFB9E;	13'h0A7C: data <= 32'hB15613FF;	13'h0A7D: data <= 32'hB18C42FE;	13'h0A7E: data <= 32'hB1C2888A;	13'h0A7F: data <= 32'hB1F8E493;	13'h0A80: data <= 32'hB22F570C;	13'h0A81: data <= 32'hB265DFE3;	13'h0A82: data <= 32'hB29C7F08;	13'h0A83: data <= 32'hB2D3346D;	13'h0A84: data <= 32'hB30A0002;	13'h0A85: data <= 32'hB340E1B6;	13'h0A86: data <= 32'hB377D97B;	13'h0A87: data <= 32'hB3AEE740;	13'h0A88: data <= 32'hB3E60AF5;	13'h0A89: data <= 32'hB41D448A;	13'h0A8A: data <= 32'hB45493F0;	13'h0A8B: data <= 32'hB48BF917;	13'h0A8C: data <= 32'hB4C373EF;	13'h0A8D: data <= 32'hB4FB0468;	13'h0A8E: data <= 32'hB532AA72;	13'h0A8F: data <= 32'hB56A65FC;	13'h0A90: data <= 32'hB5A236F8;	13'h0A91: data <= 32'hB5DA1D54;	13'h0A92: data <= 32'hB6121901;	13'h0A93: data <= 32'hB64A29EF;	13'h0A94: data <= 32'hB682500D;	13'h0A95: data <= 32'hB6BA8B4C;	13'h0A96: data <= 32'hB6F2DB9B;	13'h0A97: data <= 32'hB72B40EA;	13'h0A98: data <= 32'hB763BB29;	13'h0A99: data <= 32'hB79C4A47;	13'h0A9A: data <= 32'hB7D4EE35;	13'h0A9B: data <= 32'hB80DA6E2;	13'h0A9C: data <= 32'hB846743E;	13'h0A9D: data <= 32'hB87F5638;	13'h0A9E: data <= 32'hB8B84CC1;	13'h0A9F: data <= 32'hB8F157C7;	13'h0AA0: data <= 32'hB92A773A;	13'h0AA1: data <= 32'hB963AB0A;	13'h0AA2: data <= 32'hB99CF327;	13'h0AA3: data <= 32'hB9D64F80;	13'h0AA4: data <= 32'hBA0FC004;	13'h0AA5: data <= 32'hBA4944A3;	13'h0AA6: data <= 32'hBA82DD4D;	13'h0AA7: data <= 32'hBABC89F1;	13'h0AA8: data <= 32'hBAF64A7D;	13'h0AA9: data <= 32'hBB301EE3;	13'h0AAA: data <= 32'hBB6A0711;	13'h0AAB: data <= 32'hBBA402F6;	13'h0AAC: data <= 32'hBBDE1282;	13'h0AAD: data <= 32'hBC1835A4;	13'h0AAE: data <= 32'hBC526C4B;	13'h0AAF: data <= 32'hBC8CB667;	13'h0AB0: data <= 32'hBCC713E7;	13'h0AB1: data <= 32'hBD0184BA;	13'h0AB2: data <= 32'hBD3C08CF;	13'h0AB3: data <= 32'hBD76A016;	13'h0AB4: data <= 32'hBDB14A7D;	13'h0AB5: data <= 32'hBDEC07F4;	13'h0AB6: data <= 32'hBE26D86A;	13'h0AB7: data <= 32'hBE61BBCE;	13'h0AB8: data <= 32'hBE9CB20F;	13'h0AB9: data <= 32'hBED7BB1D;	13'h0ABA: data <= 32'hBF12D6E5;	13'h0ABB: data <= 32'hBF4E0557;	13'h0ABC: data <= 32'hBF894663;	13'h0ABD: data <= 32'hBFC499F6;	13'h0ABE: data <= 32'hC0000001;	13'h0ABF: data <= 32'hC03B7872;	13'h0AC0: data <= 32'hC0770337;	13'h0AC1: data <= 32'hC0B2A040;	13'h0AC2: data <= 32'hC0EE4F7C;	13'h0AC3: data <= 32'hC12A10D9;	13'h0AC4: data <= 32'hC165E447;	13'h0AC5: data <= 32'hC1A1C9B4;	13'h0AC6: data <= 32'hC1DDC10E;	13'h0AC7: data <= 32'hC219CA45;	13'h0AC8: data <= 32'hC255E547;	13'h0AC9: data <= 32'hC2921204;	13'h0ACA: data <= 32'hC2CE5069;	13'h0ACB: data <= 32'hC30AA066;	13'h0ACC: data <= 32'hC34701E9;	13'h0ACD: data <= 32'hC38374E1;	13'h0ACE: data <= 32'hC3BFF93C;	13'h0ACF: data <= 32'hC3FC8EE9;	13'h0AD0: data <= 32'hC43935D6;	13'h0AD1: data <= 32'hC475EDF3;	13'h0AD2: data <= 32'hC4B2B72D;	13'h0AD3: data <= 32'hC4EF9174;	13'h0AD4: data <= 32'hC52C7CB5;	13'h0AD5: data <= 32'hC56978E0;	13'h0AD6: data <= 32'hC5A685E2;	13'h0AD7: data <= 32'hC5E3A3AA;	13'h0AD8: data <= 32'hC620D227;	13'h0AD9: data <= 32'hC65E1147;	13'h0ADA: data <= 32'hC69B60F8;	13'h0ADB: data <= 32'hC6D8C129;	13'h0ADC: data <= 32'hC71631C8;	13'h0ADD: data <= 32'hC753B2C4;	13'h0ADE: data <= 32'hC791440A;	13'h0ADF: data <= 32'hC7CEE589;	13'h0AE0: data <= 32'hC80C9730;	13'h0AE1: data <= 32'hC84A58EC;	13'h0AE2: data <= 32'hC8882AAC;	13'h0AE3: data <= 32'hC8C60C5E;	13'h0AE4: data <= 32'hC903FDF0;	13'h0AE5: data <= 32'hC941FF51;	13'h0AE6: data <= 32'hC980106F;	13'h0AE7: data <= 32'hC9BE3137;	13'h0AE8: data <= 32'hC9FC6198;	13'h0AE9: data <= 32'hCA3AA180;	13'h0AEA: data <= 32'hCA78F0DE;	13'h0AEB: data <= 32'hCAB74F9F;	13'h0AEC: data <= 32'hCAF5BDB1;	13'h0AED: data <= 32'hCB343B02;	13'h0AEE: data <= 32'hCB72C781;	13'h0AEF: data <= 32'hCBB1631B;	13'h0AF0: data <= 32'hCBF00DBF;	13'h0AF1: data <= 32'hCC2EC75A;	13'h0AF2: data <= 32'hCC6D8FDB;	13'h0AF3: data <= 32'hCCAC672E;	13'h0AF4: data <= 32'hCCEB4D44;	13'h0AF5: data <= 32'hCD2A4208;	13'h0AF6: data <= 32'hCD694569;	13'h0AF7: data <= 32'hCDA85756;	13'h0AF8: data <= 32'hCDE777BB;	13'h0AF9: data <= 32'hCE26A687;	13'h0AFA: data <= 32'hCE65E3A8;	13'h0AFB: data <= 32'hCEA52F0B;	13'h0AFC: data <= 32'hCEE4889E;	13'h0AFD: data <= 32'hCF23F04F;	13'h0AFE: data <= 32'hCF63660B;	13'h0AFF: data <= 32'hCFA2E9C2;	13'h0B00: data <= 32'hCFE27B5F;	13'h0B01: data <= 32'hD0221AD2;	13'h0B02: data <= 32'hD061C807;	13'h0B03: data <= 32'hD0A182EC;	13'h0B04: data <= 32'hD0E14B70;	13'h0B05: data <= 32'hD121217F;	13'h0B06: data <= 32'hD1610507;	13'h0B07: data <= 32'hD1A0F5F7;	13'h0B08: data <= 32'hD1E0F43B;	13'h0B09: data <= 32'hD220FFC1;	13'h0B0A: data <= 32'hD2611877;	13'h0B0B: data <= 32'hD2A13E4B;	13'h0B0C: data <= 32'hD2E17129;	13'h0B0D: data <= 32'hD321B100;	13'h0B0E: data <= 32'hD361FDBD;	13'h0B0F: data <= 32'hD3A2574D;	13'h0B10: data <= 32'hD3E2BD9F;	13'h0B11: data <= 32'hD423309F;	13'h0B12: data <= 32'hD463B03B;	13'h0B13: data <= 32'hD4A43C60;	13'h0B14: data <= 32'hD4E4D4FC;	13'h0B15: data <= 32'hD52579FD;	13'h0B16: data <= 32'hD5662B4F;	13'h0B17: data <= 32'hD5A6E8E1;	13'h0B18: data <= 32'hD5E7B29F;	13'h0B19: data <= 32'hD6288876;	13'h0B1A: data <= 32'hD6696A56;	13'h0B1B: data <= 32'hD6AA5829;	13'h0B1C: data <= 32'hD6EB51DF;	13'h0B1D: data <= 32'hD72C5764;	13'h0B1E: data <= 32'hD76D68A5;	13'h0B1F: data <= 32'hD7AE8591;	13'h0B20: data <= 32'hD7EFAE13;	13'h0B21: data <= 32'hD830E21A;	13'h0B22: data <= 32'hD8722192;	13'h0B23: data <= 32'hD8B36C6A;	13'h0B24: data <= 32'hD8F4C28E;	13'h0B25: data <= 32'hD93623EA;	13'h0B26: data <= 32'hD977906E;	13'h0B27: data <= 32'hD9B90805;	13'h0B28: data <= 32'hD9FA8A9E;	13'h0B29: data <= 32'hDA3C1824;	13'h0B2A: data <= 32'hDA7DB086;	13'h0B2B: data <= 32'hDABF53B0;	13'h0B2C: data <= 32'hDB01018F;	13'h0B2D: data <= 32'hDB42BA11;	13'h0B2E: data <= 32'hDB847D23;	13'h0B2F: data <= 32'hDBC64AB2;	13'h0B30: data <= 32'hDC0822AB;	13'h0B31: data <= 32'hDC4A04FB;	13'h0B32: data <= 32'hDC8BF18E;	13'h0B33: data <= 32'hDCCDE853;	13'h0B34: data <= 32'hDD0FE937;	13'h0B35: data <= 32'hDD51F425;	13'h0B36: data <= 32'hDD94090B;	13'h0B37: data <= 32'hDDD627D7;	13'h0B38: data <= 32'hDE185075;	13'h0B39: data <= 32'hDE5A82D2;	13'h0B3A: data <= 32'hDE9CBEDB;	13'h0B3B: data <= 32'hDEDF047E;	13'h0B3C: data <= 32'hDF2153A6;	13'h0B3D: data <= 32'hDF63AC41;	13'h0B3E: data <= 32'hDFA60E3D;	13'h0B3F: data <= 32'hDFE87985;	13'h0B40: data <= 32'hE02AEE07;	13'h0B41: data <= 32'hE06D6BAF;	13'h0B42: data <= 32'hE0AFF26B;	13'h0B43: data <= 32'hE0F28228;	13'h0B44: data <= 32'hE1351AD1;	13'h0B45: data <= 32'hE177BC55;	13'h0B46: data <= 32'hE1BA66A0;	13'h0B47: data <= 32'hE1FD199E;	13'h0B48: data <= 32'hE23FD53E;	13'h0B49: data <= 32'hE282996A;	13'h0B4A: data <= 32'hE2C56611;	13'h0B4B: data <= 32'hE3083B1F;	13'h0B4C: data <= 32'hE34B1881;	13'h0B4D: data <= 32'hE38DFE23;	13'h0B4E: data <= 32'hE3D0EBF3;	13'h0B4F: data <= 32'hE413E1DD;	13'h0B50: data <= 32'hE456DFCE;	13'h0B51: data <= 32'hE499E5B2;	13'h0B52: data <= 32'hE4DCF377;	13'h0B53: data <= 32'hE5200909;	13'h0B54: data <= 32'hE5632654;	13'h0B55: data <= 32'hE5A64B47;	13'h0B56: data <= 32'hE5E977CC;	13'h0B57: data <= 32'hE62CABD1;	13'h0B58: data <= 32'hE66FE743;	13'h0B59: data <= 32'hE6B32A0E;	13'h0B5A: data <= 32'hE6F6741F;	13'h0B5B: data <= 32'hE739C563;	13'h0B5C: data <= 32'hE77D1DC6;	13'h0B5D: data <= 32'hE7C07D34;	13'h0B5E: data <= 32'hE803E39C;	13'h0B5F: data <= 32'hE84750E8;	13'h0B60: data <= 32'hE88AC506;	13'h0B61: data <= 32'hE8CE3FE2;	13'h0B62: data <= 32'hE911C16A;	13'h0B63: data <= 32'hE9554989;	13'h0B64: data <= 32'hE998D82C;	13'h0B65: data <= 32'hE9DC6D3F;	13'h0B66: data <= 32'hEA2008B0;	13'h0B67: data <= 32'hEA63AA6B;	13'h0B68: data <= 32'hEAA7525C;	13'h0B69: data <= 32'hEAEB0070;	13'h0B6A: data <= 32'hEB2EB494;	13'h0B6B: data <= 32'hEB726EB3;	13'h0B6C: data <= 32'hEBB62EBC;	13'h0B6D: data <= 32'hEBF9F499;	13'h0B6E: data <= 32'hEC3DC038;	13'h0B6F: data <= 32'hEC819185;	13'h0B70: data <= 32'hECC5686D;	13'h0B71: data <= 32'hED0944DB;	13'h0B72: data <= 32'hED4D26BE;	13'h0B73: data <= 32'hED910E00;	13'h0B74: data <= 32'hEDD4FA8F;	13'h0B75: data <= 32'hEE18EC57;	13'h0B76: data <= 32'hEE5CE345;	13'h0B77: data <= 32'hEEA0DF44;	13'h0B78: data <= 32'hEEE4E042;	13'h0B79: data <= 32'hEF28E62B;	13'h0B7A: data <= 32'hEF6CF0EB;	13'h0B7B: data <= 32'hEFB1006F;	13'h0B7C: data <= 32'hEFF514A3;	13'h0B7D: data <= 32'hF0392D74;	13'h0B7E: data <= 32'hF07D4ACE;	13'h0B7F: data <= 32'hF0C16C9D;	13'h0B80: data <= 32'hF10592CE;	13'h0B81: data <= 32'hF149BD4D;	13'h0B82: data <= 32'hF18DEC08;	13'h0B83: data <= 32'hF1D21EE9;	13'h0B84: data <= 32'hF21655DD;	13'h0B85: data <= 32'hF25A90D2;	13'h0B86: data <= 32'hF29ECFB3;	13'h0B87: data <= 32'hF2E3126D;	13'h0B88: data <= 32'hF32758EB;	13'h0B89: data <= 32'hF36BA31B;	13'h0B8A: data <= 32'hF3AFF0E9;	13'h0B8B: data <= 32'hF3F44241;	13'h0B8C: data <= 32'hF438970F;	13'h0B8D: data <= 32'hF47CEF40;	13'h0B8E: data <= 32'hF4C14AC1;	13'h0B8F: data <= 32'hF505A97C;	13'h0B90: data <= 32'hF54A0B60;	13'h0B91: data <= 32'hF58E7058;	13'h0B92: data <= 32'hF5D2D851;	13'h0B93: data <= 32'hF6174337;	13'h0B94: data <= 32'hF65BB0F5;	13'h0B95: data <= 32'hF6A0217A;	13'h0B96: data <= 32'hF6E494B0;	13'h0B97: data <= 32'hF7290A85;	13'h0B98: data <= 32'hF76D82E4;	13'h0B99: data <= 32'hF7B1FDBA;	13'h0B9A: data <= 32'hF7F67AF3;	13'h0B9B: data <= 32'hF83AFA7B;	13'h0B9C: data <= 32'hF87F7C40;	13'h0B9D: data <= 32'hF8C4002C;	13'h0B9E: data <= 32'hF908862D;	13'h0B9F: data <= 32'hF94D0E2E;	13'h0BA0: data <= 32'hF991981D;	13'h0BA1: data <= 32'hF9D623E5;	13'h0BA2: data <= 32'hFA1AB172;	13'h0BA3: data <= 32'hFA5F40B1;	13'h0BA4: data <= 32'hFAA3D18F;	13'h0BA5: data <= 32'hFAE863F7;	13'h0BA6: data <= 32'hFB2CF7D6;	13'h0BA7: data <= 32'hFB718D17;	13'h0BA8: data <= 32'hFBB623A8;	13'h0BA9: data <= 32'hFBFABB75;	13'h0BAA: data <= 32'hFC3F546A;	13'h0BAB: data <= 32'hFC83EE72;	13'h0BAC: data <= 32'hFCC8897B;	13'h0BAD: data <= 32'hFD0D2571;	13'h0BAE: data <= 32'hFD51C240;	13'h0BAF: data <= 32'hFD965FD4;	13'h0BB0: data <= 32'hFDDAFE1A;	13'h0BB1: data <= 32'hFE1F9CFE;	13'h0BB2: data <= 32'hFE643C6B;	13'h0BB3: data <= 32'hFEA8DC4F;	13'h0BB4: data <= 32'hFEED7C96;	13'h0BB5: data <= 32'hFF321D2C;	13'h0BB6: data <= 32'hFF76BDFC;	13'h0BB7: data <= 32'hFFBB5EF5;	13'h0BB8: data <= 32'h00887CBF;	13'h0BB9: data <= 32'h004B8DB2;	13'h0BBA: data <= 32'h000E9EA6;	13'h0BBB: data <= 32'hFFD1AF9B;	13'h0BBC: data <= 32'hFF94C08F;	13'h0BBD: data <= 32'hFF57D183;	13'h0BBE: data <= 32'hFF1AE277;	13'h0BBF: data <= 32'hFEDDF36B;	13'h0BC0: data <= 32'hFEA1045F;	13'h0BC1: data <= 32'hFE641553;	13'h0BC2: data <= 32'hFE272647;	13'h0BC3: data <= 32'hFDEA373B;	13'h0BC4: data <= 32'hFDAD482F;	13'h0BC5: data <= 32'hFD705923;	13'h0BC6: data <= 32'hFD336A17;	13'h0BC7: data <= 32'hFCF67B0A;	13'h0BC8: data <= 32'hFCB98BFE;	13'h0BC9: data <= 32'hFC7C9CF2;	13'h0BCA: data <= 32'hFC3FADE6;	13'h0BCB: data <= 32'hFC02BEDA;	13'h0BCC: data <= 32'hFBC5CFCE;	13'h0BCD: data <= 32'hFB88E0C2;	13'h0BCE: data <= 32'hFB4BF1B6;	13'h0BCF: data <= 32'hFB0F02AA;	13'h0BD0: data <= 32'hFAD2139E;	13'h0BD1: data <= 32'hFA952492;	13'h0BD2: data <= 32'hFA583586;	13'h0BD3: data <= 32'hFA1B467A;	13'h0BD4: data <= 32'hF9DE576E;	13'h0BD5: data <= 32'hF9A16861;	13'h0BD6: data <= 32'hF9647955;	13'h0BD7: data <= 32'hF929E31A;	13'h0BD8: data <= 32'hF8F05218;	13'h0BD9: data <= 32'hF8B6C115;	13'h0BDA: data <= 32'hF87D3013;	13'h0BDB: data <= 32'hF8439F11;	13'h0BDC: data <= 32'hF80A0E0E;	13'h0BDD: data <= 32'hF7D07D0C;	13'h0BDE: data <= 32'hF796EC0A;	13'h0BDF: data <= 32'hF75D5B07;	13'h0BE0: data <= 32'hF723CA05;	13'h0BE1: data <= 32'hF6EA3903;	13'h0BE2: data <= 32'hF6B0A800;	13'h0BE3: data <= 32'hF67716FE;	13'h0BE4: data <= 32'hF63D85FC;	13'h0BE5: data <= 32'hF603F4F9;	13'h0BE6: data <= 32'hF5CA63F7;	13'h0BE7: data <= 32'hF590D2F5;	13'h0BE8: data <= 32'hF55741F3;	13'h0BE9: data <= 32'hF51DB0F0;	13'h0BEA: data <= 32'hF4E41FEE;	13'h0BEB: data <= 32'hF4AA8EEC;	13'h0BEC: data <= 32'hF470FDE9;	13'h0BED: data <= 32'hF4376CE7;	13'h0BEE: data <= 32'hF3FDDBE5;	13'h0BEF: data <= 32'hF3C44AE2;	13'h0BF0: data <= 32'hF38AB9E0;	13'h0BF1: data <= 32'hF35128DE;	13'h0BF2: data <= 32'hF31797DB;	13'h0BF3: data <= 32'hF2DE06D9;	13'h0BF4: data <= 32'hF2A475D7;	13'h0BF5: data <= 32'hF26D3BFB;	13'h0BF6: data <= 32'hF2399BE4;	13'h0BF7: data <= 32'hF205FBCE;	13'h0BF8: data <= 32'hF1D25BB7;	13'h0BF9: data <= 32'hF19EBBA1;	13'h0BFA: data <= 32'hF16B1B8A;	13'h0BFB: data <= 32'hF1377B73;	13'h0BFC: data <= 32'hF103DB5D;	13'h0BFD: data <= 32'hF0D03B46;	13'h0BFE: data <= 32'hF09C9B30;	13'h0BFF: data <= 32'hF068FB19;	13'h0C00: data <= 32'hF0355B02;	13'h0C01: data <= 32'hF001BAEC;	13'h0C02: data <= 32'hEFCE1AD5;	13'h0C03: data <= 32'hEF9A7ABF;	13'h0C04: data <= 32'hEF66DAA8;	13'h0C05: data <= 32'hEF333A91;	13'h0C06: data <= 32'hEEFF9A7B;	13'h0C07: data <= 32'hEECBFA64;	13'h0C08: data <= 32'hEE985A4E;	13'h0C09: data <= 32'hEE64BA37;	13'h0C0A: data <= 32'hEE311A20;	13'h0C0B: data <= 32'hEDFD7A0A;	13'h0C0C: data <= 32'hEDC9D9F3;	13'h0C0D: data <= 32'hED9639DD;	13'h0C0E: data <= 32'hED6299C6;	13'h0C0F: data <= 32'hED2EF9AF;	13'h0C10: data <= 32'hECFB5999;	13'h0C11: data <= 32'hECC7B982;	13'h0C12: data <= 32'hEC94196C;	13'h0C13: data <= 32'hEC613882;	13'h0C14: data <= 32'hEC35CF5B;	13'h0C15: data <= 32'hEC0A6633;	13'h0C16: data <= 32'hEBDEFD0C;	13'h0C17: data <= 32'hEBB393E4;	13'h0C18: data <= 32'hEB882ABC;	13'h0C19: data <= 32'hEB5CC195;	13'h0C1A: data <= 32'hEB31586D;	13'h0C1B: data <= 32'hEB05EF46;	13'h0C1C: data <= 32'hEADA861E;	13'h0C1D: data <= 32'hEAAF1CF7;	13'h0C1E: data <= 32'hEA83B3CF;	13'h0C1F: data <= 32'hEA584AA8;	13'h0C20: data <= 32'hEA2CE180;	13'h0C21: data <= 32'hEA017859;	13'h0C22: data <= 32'hE9D60F31;	13'h0C23: data <= 32'hE9AAA60A;	13'h0C24: data <= 32'hE97F3CE2;	13'h0C25: data <= 32'hE953D3BB;	13'h0C26: data <= 32'hE9286A93;	13'h0C27: data <= 32'hE8FD016C;	13'h0C28: data <= 32'hE8D19844;	13'h0C29: data <= 32'hE8A62F1D;	13'h0C2A: data <= 32'hE87AC5F5;	13'h0C2B: data <= 32'hE84F5CCE;	13'h0C2C: data <= 32'hE823F3A6;	13'h0C2D: data <= 32'hE7F88A7F;	13'h0C2E: data <= 32'hE7CD2157;	13'h0C2F: data <= 32'hE7A1B830;	13'h0C30: data <= 32'hE7764F08;	13'h0C31: data <= 32'hE74AE5E0;	13'h0C32: data <= 32'hE726A6F2;	13'h0C33: data <= 32'hE70455D8;	13'h0C34: data <= 32'hE6E204BE;	13'h0C35: data <= 32'hE6BFB3A3;	13'h0C36: data <= 32'hE69D6289;	13'h0C37: data <= 32'hE67B116F;	13'h0C38: data <= 32'hE658C055;	13'h0C39: data <= 32'hE6366F3B;	13'h0C3A: data <= 32'hE6141E20;	13'h0C3B: data <= 32'hE5F1CD06;	13'h0C3C: data <= 32'hE5CF7BEC;	13'h0C3D: data <= 32'hE5AD2AD2;	13'h0C3E: data <= 32'hE58AD9B8;	13'h0C3F: data <= 32'hE568889D;	13'h0C40: data <= 32'hE5463783;	13'h0C41: data <= 32'hE523E669;	13'h0C42: data <= 32'hE501954F;	13'h0C43: data <= 32'hE4DF4435;	13'h0C44: data <= 32'hE4BCF31A;	13'h0C45: data <= 32'hE49AA200;	13'h0C46: data <= 32'hE47850E6;	13'h0C47: data <= 32'hE455FFCC;	13'h0C48: data <= 32'hE433AEB2;	13'h0C49: data <= 32'hE4115D97;	13'h0C4A: data <= 32'hE3EF0C7D;	13'h0C4B: data <= 32'hE3CCBB63;	13'h0C4C: data <= 32'hE3AA6A49;	13'h0C4D: data <= 32'hE388192F;	13'h0C4E: data <= 32'hE365C814;	13'h0C4F: data <= 32'hE34376FA;	13'h0C50: data <= 32'hE324C44E;	13'h0C51: data <= 32'hE309E9F6;	13'h0C52: data <= 32'hE2EF0F9E;	13'h0C53: data <= 32'hE2D43547;	13'h0C54: data <= 32'hE2B95AEF;	13'h0C55: data <= 32'hE29E8097;	13'h0C56: data <= 32'hE283A640;	13'h0C57: data <= 32'hE268CBE8;	13'h0C58: data <= 32'hE24DF190;	13'h0C59: data <= 32'hE2331739;	13'h0C5A: data <= 32'hE2183CE1;	13'h0C5B: data <= 32'hE1FD6289;	13'h0C5C: data <= 32'hE1E28832;	13'h0C5D: data <= 32'hE1C7ADDA;	13'h0C5E: data <= 32'hE1ACD382;	13'h0C5F: data <= 32'hE191F92A;	13'h0C60: data <= 32'hE1771ED3;	13'h0C61: data <= 32'hE15C447B;	13'h0C62: data <= 32'hE1416A23;	13'h0C63: data <= 32'hE1268FCC;	13'h0C64: data <= 32'hE10BB574;	13'h0C65: data <= 32'hE0F0DB1C;	13'h0C66: data <= 32'hE0D600C5;	13'h0C67: data <= 32'hE0BB266D;	13'h0C68: data <= 32'hE0A04C15;	13'h0C69: data <= 32'hE08571BE;	13'h0C6A: data <= 32'hE06A9766;	13'h0C6B: data <= 32'hE04FBD0E;	13'h0C6C: data <= 32'hE034E2B6;	13'h0C6D: data <= 32'hE01A085F;	13'h0C6E: data <= 32'hDFFFF5B0;	13'h0C6F: data <= 32'hDFE9657C;	13'h0C70: data <= 32'hDFD2D548;	13'h0C71: data <= 32'hDFBC4513;	13'h0C72: data <= 32'hDFA5B4DF;	13'h0C73: data <= 32'hDF8F24AA;	13'h0C74: data <= 32'hDF789476;	13'h0C75: data <= 32'hDF620441;	13'h0C76: data <= 32'hDF4B740D;	13'h0C77: data <= 32'hDF34E3D9;	13'h0C78: data <= 32'hDF1E53A4;	13'h0C79: data <= 32'hDF07C370;	13'h0C7A: data <= 32'hDEF1333B;	13'h0C7B: data <= 32'hDEDAA307;	13'h0C7C: data <= 32'hDEC412D3;	13'h0C7D: data <= 32'hDEAD829E;	13'h0C7E: data <= 32'hDE96F26A;	13'h0C7F: data <= 32'hDE806235;	13'h0C80: data <= 32'hDE69D201;	13'h0C81: data <= 32'hDE5341CC;	13'h0C82: data <= 32'hDE3CB198;	13'h0C83: data <= 32'hDE262164;	13'h0C84: data <= 32'hDE0F912F;	13'h0C85: data <= 32'hDDF900FB;	13'h0C86: data <= 32'hDDE270C6;	13'h0C87: data <= 32'hDDCBE092;	13'h0C88: data <= 32'hDDB5505E;	13'h0C89: data <= 32'hDD9EC029;	13'h0C8A: data <= 32'hDD882FF5;	13'h0C8B: data <= 32'hDD719FC0;	13'h0C8C: data <= 32'hDD5B0F8C;	13'h0C8D: data <= 32'hDD44FCCC;	13'h0C8E: data <= 32'hDD2EFB59;	13'h0C8F: data <= 32'hDD18F9E7;	13'h0C90: data <= 32'hDD02F874;	13'h0C91: data <= 32'hDCECF702;	13'h0C92: data <= 32'hDCD6F590;	13'h0C93: data <= 32'hDCC0F41D;	13'h0C94: data <= 32'hDCAAF2AB;	13'h0C95: data <= 32'hDC94F138;	13'h0C96: data <= 32'hDC7EEFC6;	13'h0C97: data <= 32'hDC68EE54;	13'h0C98: data <= 32'hDC52ECE1;	13'h0C99: data <= 32'hDC3CEB6F;	13'h0C9A: data <= 32'hDC26E9FC;	13'h0C9B: data <= 32'hDC10E88A;	13'h0C9C: data <= 32'hDBFAE718;	13'h0C9D: data <= 32'hDBE4E5A5;	13'h0C9E: data <= 32'hDBCEE433;	13'h0C9F: data <= 32'hDBB8E2C0;	13'h0CA0: data <= 32'hDBA2E14E;	13'h0CA1: data <= 32'hDB8CDFDC;	13'h0CA2: data <= 32'hDB76DE69;	13'h0CA3: data <= 32'hDB60DCF7;	13'h0CA4: data <= 32'hDB4ADB84;	13'h0CA5: data <= 32'hDB34DA12;	13'h0CA6: data <= 32'hDB1ED8A0;	13'h0CA7: data <= 32'hDB08D72D;	13'h0CA8: data <= 32'hDAF2D5BB;	13'h0CA9: data <= 32'hDADCD448;	13'h0CAA: data <= 32'hDAC6D2D6;	13'h0CAB: data <= 32'hDAAF3342;	13'h0CAC: data <= 32'hDA966288;	13'h0CAD: data <= 32'hDA7D91CE;	13'h0CAE: data <= 32'hDA64C114;	13'h0CAF: data <= 32'hDA4BF05A;	13'h0CB0: data <= 32'hDA331F9F;	13'h0CB1: data <= 32'hDA1A4EE5;	13'h0CB2: data <= 32'hDA017E2B;	13'h0CB3: data <= 32'hD9E8AD71;	13'h0CB4: data <= 32'hD9CFDCB7;	13'h0CB5: data <= 32'hD9B70BFD;	13'h0CB6: data <= 32'hD99E3B43;	13'h0CB7: data <= 32'hD9856A89;	13'h0CB8: data <= 32'hD96C99CF;	13'h0CB9: data <= 32'hD953C914;	13'h0CBA: data <= 32'hD93AF85A;	13'h0CBB: data <= 32'hD92227A0;	13'h0CBC: data <= 32'hD90956E6;	13'h0CBD: data <= 32'hD8F0862C;	13'h0CBE: data <= 32'hD8D7B572;	13'h0CBF: data <= 32'hD8BEE4B8;	13'h0CC0: data <= 32'hD8A613FE;	13'h0CC1: data <= 32'hD88D4344;	13'h0CC2: data <= 32'hD8747289;	13'h0CC3: data <= 32'hD85BA1CF;	13'h0CC4: data <= 32'hD842D115;	13'h0CC5: data <= 32'hD82A005B;	13'h0CC6: data <= 32'hD8112FA1;	13'h0CC7: data <= 32'hD7F85EE7;	13'h0CC8: data <= 32'hD7DF8E2D;	13'h0CC9: data <= 32'hD7C54297;	13'h0CCA: data <= 32'hD7A704B8;	13'h0CCB: data <= 32'hD788C6D9;	13'h0CCC: data <= 32'hD76A88FA;	13'h0CCD: data <= 32'hD74C4B1B;	13'h0CCE: data <= 32'hD72E0D3C;	13'h0CCF: data <= 32'hD70FCF5D;	13'h0CD0: data <= 32'hD6F1917E;	13'h0CD1: data <= 32'hD6D3539E;	13'h0CD2: data <= 32'hD6B515BF;	13'h0CD3: data <= 32'hD696D7E0;	13'h0CD4: data <= 32'hD6789A01;	13'h0CD5: data <= 32'hD65A5C22;	13'h0CD6: data <= 32'hD63C1E43;	13'h0CD7: data <= 32'hD61DE064;	13'h0CD8: data <= 32'hD5FFA285;	13'h0CD9: data <= 32'hD5E164A6;	13'h0CDA: data <= 32'hD5C326C7;	13'h0CDB: data <= 32'hD5A4E8E8;	13'h0CDC: data <= 32'hD586AB09;	13'h0CDD: data <= 32'hD5686D29;	13'h0CDE: data <= 32'hD54A2F4A;	13'h0CDF: data <= 32'hD52BF16B;	13'h0CE0: data <= 32'hD50DB38C;	13'h0CE1: data <= 32'hD4EF75AD;	13'h0CE2: data <= 32'hD4D137CE;	13'h0CE3: data <= 32'hD4B2F9EF;	13'h0CE4: data <= 32'hD494BC10;	13'h0CE5: data <= 32'hD4767E31;	13'h0CE6: data <= 32'hD4584052;	13'h0CE7: data <= 32'hD43A0273;	13'h0CE8: data <= 32'hD4154765;	13'h0CE9: data <= 32'hD3F0586D;	13'h0CEA: data <= 32'hD3CB6976;	13'h0CEB: data <= 32'hD3A67A7F;	13'h0CEC: data <= 32'hD3818B87;	13'h0CED: data <= 32'hD35C9C90;	13'h0CEE: data <= 32'hD337AD98;	13'h0CEF: data <= 32'hD312BEA1;	13'h0CF0: data <= 32'hD2EDCFAA;	13'h0CF1: data <= 32'hD2C8E0B2;	13'h0CF2: data <= 32'hD2A3F1BB;	13'h0CF3: data <= 32'hD27F02C3;	13'h0CF4: data <= 32'hD25A13CC;	13'h0CF5: data <= 32'hD23524D5;	13'h0CF6: data <= 32'hD21035DD;	13'h0CF7: data <= 32'hD1EB46E6;	13'h0CF8: data <= 32'hD1C657EE;	13'h0CF9: data <= 32'hD1A168F7;	13'h0CFA: data <= 32'hD17C7A00;	13'h0CFB: data <= 32'hD1578B08;	13'h0CFC: data <= 32'hD1329C11;	13'h0CFD: data <= 32'hD10DAD19;	13'h0CFE: data <= 32'hD0E8BE22;	13'h0CFF: data <= 32'hD0C3CF2B;	13'h0D00: data <= 32'hD09EE033;	13'h0D01: data <= 32'hD079F13C;	13'h0D02: data <= 32'hD0550244;	13'h0D03: data <= 32'hD030134D;	13'h0D04: data <= 32'hD00B2456;	13'h0D05: data <= 32'hCFE6355E;	13'h0D06: data <= 32'hCFBCA46A;	13'h0D07: data <= 32'hCF90C277;	13'h0D08: data <= 32'hCF64E084;	13'h0D09: data <= 32'hCF38FE90;	13'h0D0A: data <= 32'hCF0D1C9D;	13'h0D0B: data <= 32'hCEE13AAA;	13'h0D0C: data <= 32'hCEB558B7;	13'h0D0D: data <= 32'hCE8976C4;	13'h0D0E: data <= 32'hCE5D94D1;	13'h0D0F: data <= 32'hCE31B2DE;	13'h0D10: data <= 32'hCE05D0EB;	13'h0D11: data <= 32'hCDD9EEF8;	13'h0D12: data <= 32'hCDAE0D05;	13'h0D13: data <= 32'hCD822B12;	13'h0D14: data <= 32'hCD56491E;	13'h0D15: data <= 32'hCD2A672B;	13'h0D16: data <= 32'hCCFE8538;	13'h0D17: data <= 32'hCCD2A345;	13'h0D18: data <= 32'hCCA6C152;	13'h0D19: data <= 32'hCC7ADF5F;	13'h0D1A: data <= 32'hCC4EFD6C;	13'h0D1B: data <= 32'hCC231B79;	13'h0D1C: data <= 32'hCBF73986;	13'h0D1D: data <= 32'hCBCB5793;	13'h0D1E: data <= 32'hCB9F759F;	13'h0D1F: data <= 32'hCB7393AC;	13'h0D20: data <= 32'hCB47B1B9;	13'h0D21: data <= 32'hCB1BCFC6;	13'h0D22: data <= 32'hCAEFEDD3;	13'h0D23: data <= 32'hCAC40BE0;	13'h0D24: data <= 32'hCA95CAF4;	13'h0D25: data <= 32'hCA6363D6;	13'h0D26: data <= 32'hCA30FCB8;	13'h0D27: data <= 32'hC9FE9599;	13'h0D28: data <= 32'hC9CC2E7B;	13'h0D29: data <= 32'hC999C75C;	13'h0D2A: data <= 32'hC967603E;	13'h0D2B: data <= 32'hC934F91F;	13'h0D2C: data <= 32'hC9029201;	13'h0D2D: data <= 32'hC8D02AE2;	13'h0D2E: data <= 32'hC89DC3C4;	13'h0D2F: data <= 32'hC86B5CA5;	13'h0D30: data <= 32'hC838F587;	13'h0D31: data <= 32'hC8068E68;	13'h0D32: data <= 32'hC7D4274A;	13'h0D33: data <= 32'hC7A1C02C;	13'h0D34: data <= 32'hC76F590D;	13'h0D35: data <= 32'hC73CF1EF;	13'h0D36: data <= 32'hC70A8AD0;	13'h0D37: data <= 32'hC6D823B2;	13'h0D38: data <= 32'hC6A5BC93;	13'h0D39: data <= 32'hC6735575;	13'h0D3A: data <= 32'hC640EE56;	13'h0D3B: data <= 32'hC60E8738;	13'h0D3C: data <= 32'hC5DC2019;	13'h0D3D: data <= 32'hC5A9B8FB;	13'h0D3E: data <= 32'hC57751DC;	13'h0D3F: data <= 32'hC544EABE;	13'h0D40: data <= 32'hC51283A0;	13'h0D41: data <= 32'hC4E01C81;	13'h0D42: data <= 32'hC4AD7081;	13'h0D43: data <= 32'hC47698D0;	13'h0D44: data <= 32'hC43FC11E;	13'h0D45: data <= 32'hC408E96D;	13'h0D46: data <= 32'hC3D211BC;	13'h0D47: data <= 32'hC39B3A0B;	13'h0D48: data <= 32'hC364625A;	13'h0D49: data <= 32'hC32D8AA9;	13'h0D4A: data <= 32'hC2F6B2F8;	13'h0D4B: data <= 32'hC2BFDB47;	13'h0D4C: data <= 32'hC2890396;	13'h0D4D: data <= 32'hC2522BE5;	13'h0D4E: data <= 32'hC21B5434;	13'h0D4F: data <= 32'hC1E47C83;	13'h0D50: data <= 32'hC1ADA4D2;	13'h0D51: data <= 32'hC176CD21;	13'h0D52: data <= 32'hC13FF570;	13'h0D53: data <= 32'hC1091DBF;	13'h0D54: data <= 32'hC0D2460E;	13'h0D55: data <= 32'hC09B6E5D;	13'h0D56: data <= 32'hC06496AC;	13'h0D57: data <= 32'hC02DBEFB;	13'h0D58: data <= 32'hBFF6E74A;	13'h0D59: data <= 32'hBFC00F99;	13'h0D5A: data <= 32'hBF8937E8;	13'h0D5B: data <= 32'hBF526036;	13'h0D5C: data <= 32'hBF1B8885;	13'h0D5D: data <= 32'hBEE4B0D4;	13'h0D5E: data <= 32'hBEADD923;	13'h0D5F: data <= 32'hBE770172;	13'h0D60: data <= 32'hBE4029C1;	13'h0D61: data <= 32'hBE08C4A3;	13'h0D62: data <= 32'hBDD13243;	13'h0D63: data <= 32'hBD999FE3;	13'h0D64: data <= 32'hBD620D83;	13'h0D65: data <= 32'hBD2A7B23;	13'h0D66: data <= 32'hBCF2E8C3;	13'h0D67: data <= 32'hBCBB5663;	13'h0D68: data <= 32'hBC83C403;	13'h0D69: data <= 32'hBC4C31A3;	13'h0D6A: data <= 32'hBC149F43;	13'h0D6B: data <= 32'hBBDD0CE3;	13'h0D6C: data <= 32'hBBA57A83;	13'h0D6D: data <= 32'hBB6DE823;	13'h0D6E: data <= 32'hBB3655C3;	13'h0D6F: data <= 32'hBAFEC363;	13'h0D70: data <= 32'hBAC73103;	13'h0D71: data <= 32'hBA8F9EA3;	13'h0D72: data <= 32'hBA580C43;	13'h0D73: data <= 32'hBA2079E3;	13'h0D74: data <= 32'hB9E8E783;	13'h0D75: data <= 32'hB9B15523;	13'h0D76: data <= 32'hB979C2C3;	13'h0D77: data <= 32'hB9423063;	13'h0D78: data <= 32'hB90A9E03;	13'h0D79: data <= 32'hB8D30BA3;	13'h0D7A: data <= 32'hB89B7943;	13'h0D7B: data <= 32'hB863E6E3;	13'h0D7C: data <= 32'hB82C5483;	13'h0D7D: data <= 32'hB7F4C223;	13'h0D7E: data <= 32'hB7BD2FC3;	13'h0D7F: data <= 32'hB7871141;	13'h0D80: data <= 32'hB752B0FE;	13'h0D81: data <= 32'hB71E50BB;	13'h0D82: data <= 32'hB6E9F078;	13'h0D83: data <= 32'hB6B59035;	13'h0D84: data <= 32'hB6812FF2;	13'h0D85: data <= 32'hB64CCFAE;	13'h0D86: data <= 32'hB6186F6B;	13'h0D87: data <= 32'hB5E40F28;	13'h0D88: data <= 32'hB5AFAEE5;	13'h0D89: data <= 32'hB57B4EA2;	13'h0D8A: data <= 32'hB546EE5F;	13'h0D8B: data <= 32'hB5128E1B;	13'h0D8C: data <= 32'hB4DE2DD8;	13'h0D8D: data <= 32'hB4A9CD95;	13'h0D8E: data <= 32'hB4756D52;	13'h0D8F: data <= 32'hB4410D0F;	13'h0D90: data <= 32'hB40CACCC;	13'h0D91: data <= 32'hB3D84C88;	13'h0D92: data <= 32'hB3A3EC45;	13'h0D93: data <= 32'hB36F8C02;	13'h0D94: data <= 32'hB33B2BBF;	13'h0D95: data <= 32'hB306CB7C;	13'h0D96: data <= 32'hB2D26B39;	13'h0D97: data <= 32'hB29E0AF5;	13'h0D98: data <= 32'hB269AAB2;	13'h0D99: data <= 32'hB2354A6F;	13'h0D9A: data <= 32'hB200EA2C;	13'h0D9B: data <= 32'hB1CC89E9;	13'h0D9C: data <= 32'hB19829A6;	13'h0D9D: data <= 32'hB164B5A7;	13'h0D9E: data <= 32'hB1366CBE;	13'h0D9F: data <= 32'hB10823D6;	13'h0DA0: data <= 32'hB0D9DAEE;	13'h0DA1: data <= 32'hB0AB9206;	13'h0DA2: data <= 32'hB07D491E;	13'h0DA3: data <= 32'hB04F0036;	13'h0DA4: data <= 32'hB020B74E;	13'h0DA5: data <= 32'hAFF26E66;	13'h0DA6: data <= 32'hAFC4257E;	13'h0DA7: data <= 32'hAF95DC96;	13'h0DA8: data <= 32'hAF6793AD;	13'h0DA9: data <= 32'hAF394AC5;	13'h0DAA: data <= 32'hAF0B01DD;	13'h0DAB: data <= 32'hAEDCB8F5;	13'h0DAC: data <= 32'hAEAE700D;	13'h0DAD: data <= 32'hAE802725;	13'h0DAE: data <= 32'hAE51DE3D;	13'h0DAF: data <= 32'hAE239555;	13'h0DB0: data <= 32'hADF54C6D;	13'h0DB1: data <= 32'hADC70384;	13'h0DB2: data <= 32'hAD98BA9C;	13'h0DB3: data <= 32'hAD6A71B4;	13'h0DB4: data <= 32'hAD3C28CC;	13'h0DB5: data <= 32'hAD0DDFE4;	13'h0DB6: data <= 32'hACDF96FC;	13'h0DB7: data <= 32'hACB14E14;	13'h0DB8: data <= 32'hAC83052C;	13'h0DB9: data <= 32'hAC54BC44;	13'h0DBA: data <= 32'hAC26735C;	13'h0DBB: data <= 32'hABF82A73;	13'h0DBC: data <= 32'hABD0F5CE;	13'h0DBD: data <= 32'hABAB04C7;	13'h0DBE: data <= 32'hAB8513BF;	13'h0DBF: data <= 32'hAB5F22B8;	13'h0DC0: data <= 32'hAB3931B0;	13'h0DC1: data <= 32'hAB1340A9;	13'h0DC2: data <= 32'hAAED4FA2;	13'h0DC3: data <= 32'hAAC75E9A;	13'h0DC4: data <= 32'hAAA16D93;	13'h0DC5: data <= 32'hAA7B7C8B;	13'h0DC6: data <= 32'hAA558B84;	13'h0DC7: data <= 32'hAA2F9A7D;	13'h0DC8: data <= 32'hAA09A975;	13'h0DC9: data <= 32'hA9E3B86E;	13'h0DCA: data <= 32'hA9BDC767;	13'h0DCB: data <= 32'hA997D65F;	13'h0DCC: data <= 32'hA971E558;	13'h0DCD: data <= 32'hA94BF450;	13'h0DCE: data <= 32'hA9260349;	13'h0DCF: data <= 32'hA9001242;	13'h0DD0: data <= 32'hA8DA213A;	13'h0DD1: data <= 32'hA8B43033;	13'h0DD2: data <= 32'hA88E3F2C;	13'h0DD3: data <= 32'hA8684E24;	13'h0DD4: data <= 32'hA8425D1D;	13'h0DD5: data <= 32'hA81C6C15;	13'h0DD6: data <= 32'hA7F67B0E;	13'h0DD7: data <= 32'hA7D08A07;	13'h0DD8: data <= 32'hA7AA98FF;	13'h0DD9: data <= 32'hA784A7F8;	13'h0DDA: data <= 32'hA7647572;	13'h0DDB: data <= 32'hA7490C58;	13'h0DDC: data <= 32'hA72DA33F;	13'h0DDD: data <= 32'hA7123A25;	13'h0DDE: data <= 32'hA6F6D10B;	13'h0DDF: data <= 32'hA6DB67F2;	13'h0DE0: data <= 32'hA6BFFED8;	13'h0DE1: data <= 32'hA6A495BE;	13'h0DE2: data <= 32'hA6892CA4;	13'h0DE3: data <= 32'hA66DC38B;	13'h0DE4: data <= 32'hA6525A71;	13'h0DE5: data <= 32'hA636F157;	13'h0DE6: data <= 32'hA61B883E;	13'h0DE7: data <= 32'hA6001F24;	13'h0DE8: data <= 32'hA5E4B60A;	13'h0DE9: data <= 32'hA5C94CF1;	13'h0DEA: data <= 32'hA5ADE3D7;	13'h0DEB: data <= 32'hA5927ABD;	13'h0DEC: data <= 32'hA57711A3;	13'h0DED: data <= 32'hA55BA88A;	13'h0DEE: data <= 32'hA5403F70;	13'h0DEF: data <= 32'hA524D656;	13'h0DF0: data <= 32'hA5096D3D;	13'h0DF1: data <= 32'hA4EE0423;	13'h0DF2: data <= 32'hA4D29B09;	13'h0DF3: data <= 32'hA4B731F0;	13'h0DF4: data <= 32'hA49BC8D6;	13'h0DF5: data <= 32'hA4805FBC;	13'h0DF6: data <= 32'hA464F6A2;	13'h0DF7: data <= 32'hA4498D89;	13'h0DF8: data <= 32'hA430EB3A;	13'h0DF9: data <= 32'hA420F628;	13'h0DFA: data <= 32'hA4110115;	13'h0DFB: data <= 32'hA4010C03;	13'h0DFC: data <= 32'hA3F116F0;	13'h0DFD: data <= 32'hA3E121DE;	13'h0DFE: data <= 32'hA3D12CCB;	13'h0DFF: data <= 32'hA3C137B8;	13'h0E00: data <= 32'hA3B142A6;	13'h0E01: data <= 32'hA3A14D93;	13'h0E02: data <= 32'hA3915881;	13'h0E03: data <= 32'hA381636E;	13'h0E04: data <= 32'hA3716E5B;	13'h0E05: data <= 32'hA3617949;	13'h0E06: data <= 32'hA3518436;	13'h0E07: data <= 32'hA3418F24;	13'h0E08: data <= 32'hA3319A11;	13'h0E09: data <= 32'hA321A4FF;	13'h0E0A: data <= 32'hA311AFEC;	13'h0E0B: data <= 32'hA301BAD9;	13'h0E0C: data <= 32'hA2F1C5C7;	13'h0E0D: data <= 32'hA2E1D0B4;	13'h0E0E: data <= 32'hA2D1DBA2;	13'h0E0F: data <= 32'hA2C1E68F;	13'h0E10: data <= 32'hA2B1F17C;	13'h0E11: data <= 32'hA2A1FC6A;	13'h0E12: data <= 32'hA2920757;	13'h0E13: data <= 32'hA2821245;	13'h0E14: data <= 32'hA2721D32;	13'h0E15: data <= 32'hA2622820;	13'h0E16: data <= 32'hA252330D;	13'h0E17: data <= 32'hA24BE49F;	13'h0E18: data <= 32'hA2463597;	13'h0E19: data <= 32'hA240868F;	13'h0E1A: data <= 32'hA23AD786;	13'h0E1B: data <= 32'hA235287E;	13'h0E1C: data <= 32'hA22F7976;	13'h0E1D: data <= 32'hA229CA6D;	13'h0E1E: data <= 32'hA2241B65;	13'h0E1F: data <= 32'hA21E6C5D;	13'h0E20: data <= 32'hA218BD54;	13'h0E21: data <= 32'hA2130E4C;	13'h0E22: data <= 32'hA20D5F44;	13'h0E23: data <= 32'hA207B03B;	13'h0E24: data <= 32'hA2020133;	13'h0E25: data <= 32'hA1FC522B;	13'h0E26: data <= 32'hA1F6A322;	13'h0E27: data <= 32'hA1F0F41A;	13'h0E28: data <= 32'hA1EB4512;	13'h0E29: data <= 32'hA1E59609;	13'h0E2A: data <= 32'hA1DFE701;	13'h0E2B: data <= 32'hA1DA37F9;	13'h0E2C: data <= 32'hA1D488F0;	13'h0E2D: data <= 32'hA1CED9E8;	13'h0E2E: data <= 32'hA1C92AE0;	13'h0E2F: data <= 32'hA1C37BD7;	13'h0E30: data <= 32'hA1BDCCCF;	13'h0E31: data <= 32'hA1B81DC7;	13'h0E32: data <= 32'hA1B26EBE;	13'h0E33: data <= 32'hA1ACBFB6;	13'h0E34: data <= 32'hA1A710AE;	13'h0E35: data <= 32'hA1A6836B;	13'h0E36: data <= 32'hA1A8E4E3;	13'h0E37: data <= 32'hA1AB465A;	13'h0E38: data <= 32'hA1ADA7D1;	13'h0E39: data <= 32'hA1B00949;	13'h0E3A: data <= 32'hA1B26AC0;	13'h0E3B: data <= 32'hA1B4CC38;	13'h0E3C: data <= 32'hA1B72DAF;	13'h0E3D: data <= 32'hA1B98F26;	13'h0E3E: data <= 32'hA1BBF09E;	13'h0E3F: data <= 32'hA1BE5215;	13'h0E40: data <= 32'hA1C0B38D;	13'h0E41: data <= 32'hA1C31504;	13'h0E42: data <= 32'hA1C5767B;	13'h0E43: data <= 32'hA1C7D7F3;	13'h0E44: data <= 32'hA1CA396A;	13'h0E45: data <= 32'hA1CC9AE2;	13'h0E46: data <= 32'hA1CEFC59;	13'h0E47: data <= 32'hA1D15DD0;	13'h0E48: data <= 32'hA1D3BF48;	13'h0E49: data <= 32'hA1D620BF;	13'h0E4A: data <= 32'hA1D88237;	13'h0E4B: data <= 32'hA1DAE3AE;	13'h0E4C: data <= 32'hA1DD4525;	13'h0E4D: data <= 32'hA1DFA69D;	13'h0E4E: data <= 32'hA1E20814;	13'h0E4F: data <= 32'hA1E4698C;	13'h0E50: data <= 32'hA1E6CB03;	13'h0E51: data <= 32'hA1E92C7A;	13'h0E52: data <= 32'hA1EB8DF2;	13'h0E53: data <= 32'hA1F00EFD;	13'h0E54: data <= 32'hA1F8CF31;	13'h0E55: data <= 32'hA2018F64;	13'h0E56: data <= 32'hA20A4F98;	13'h0E57: data <= 32'hA2130FCB;	13'h0E58: data <= 32'hA21BCFFF;	13'h0E59: data <= 32'hA2249032;	13'h0E5A: data <= 32'hA22D5066;	13'h0E5B: data <= 32'hA2361099;	13'h0E5C: data <= 32'hA23ED0CD;	13'h0E5D: data <= 32'hA2479100;	13'h0E5E: data <= 32'hA2505134;	13'h0E5F: data <= 32'hA2591167;	13'h0E60: data <= 32'hA261D19B;	13'h0E61: data <= 32'hA26A91CE;	13'h0E62: data <= 32'hA2735202;	13'h0E63: data <= 32'hA27C1235;	13'h0E64: data <= 32'hA284D269;	13'h0E65: data <= 32'hA28D929C;	13'h0E66: data <= 32'hA29652D0;	13'h0E67: data <= 32'hA29F1303;	13'h0E68: data <= 32'hA2A7D337;	13'h0E69: data <= 32'hA2B0936A;	13'h0E6A: data <= 32'hA2B9539E;	13'h0E6B: data <= 32'hA2C213D1;	13'h0E6C: data <= 32'hA2CAD405;	13'h0E6D: data <= 32'hA2D39438;	13'h0E6E: data <= 32'hA2DC546C;	13'h0E6F: data <= 32'hA2E5149F;	13'h0E70: data <= 32'hA2EDD4D3;	13'h0E71: data <= 32'hA2F6B7F7;	13'h0E72: data <= 32'hA303F936;	13'h0E73: data <= 32'hA3113A75;	13'h0E74: data <= 32'hA31E7BB4;	13'h0E75: data <= 32'hA32BBCF3;	13'h0E76: data <= 32'hA338FE31;	13'h0E77: data <= 32'hA3463F70;	13'h0E78: data <= 32'hA35380AF;	13'h0E79: data <= 32'hA360C1EE;	13'h0E7A: data <= 32'hA36E032D;	13'h0E7B: data <= 32'hA37B446C;	13'h0E7C: data <= 32'hA38885AB;	13'h0E7D: data <= 32'hA395C6EA;	13'h0E7E: data <= 32'hA3A30829;	13'h0E7F: data <= 32'hA3B04968;	13'h0E80: data <= 32'hA3BD8AA7;	13'h0E81: data <= 32'hA3CACBE5;	13'h0E82: data <= 32'hA3D80D24;	13'h0E83: data <= 32'hA3E54E63;	13'h0E84: data <= 32'hA3F28FA2;	13'h0E85: data <= 32'hA3FFD0E1;	13'h0E86: data <= 32'hA40D1220;	13'h0E87: data <= 32'hA41A535F;	13'h0E88: data <= 32'hA427949E;	13'h0E89: data <= 32'hA434D5DD;	13'h0E8A: data <= 32'hA442171C;	13'h0E8B: data <= 32'hA44F585B;	13'h0E8C: data <= 32'hA45C999A;	13'h0E8D: data <= 32'hA469DAD8;	13'h0E8E: data <= 32'hA4771C17;	13'h0E8F: data <= 32'hA4845D56;	13'h0E90: data <= 32'hA49315F2;	13'h0E91: data <= 32'hA4A25B51;	13'h0E92: data <= 32'hA4B1A0B0;	13'h0E93: data <= 32'hA4C0E60F;	13'h0E94: data <= 32'hA4D02B6E;	13'h0E95: data <= 32'hA4DF70CC;	13'h0E96: data <= 32'hA4EEB62B;	13'h0E97: data <= 32'hA4FDFB8A;	13'h0E98: data <= 32'hA50D40E9;	13'h0E99: data <= 32'hA51C8648;	13'h0E9A: data <= 32'hA52BCBA7;	13'h0E9B: data <= 32'hA53B1106;	13'h0E9C: data <= 32'hA54A5664;	13'h0E9D: data <= 32'hA5599BC3;	13'h0E9E: data <= 32'hA568E122;	13'h0E9F: data <= 32'hA5782681;	13'h0EA0: data <= 32'hA5876BE0;	13'h0EA1: data <= 32'hA596B13F;	13'h0EA2: data <= 32'hA5A5F69E;	13'h0EA3: data <= 32'hA5B53BFC;	13'h0EA4: data <= 32'hA5C4815B;	13'h0EA5: data <= 32'hA5D3C6BA;	13'h0EA6: data <= 32'hA5E30C19;	13'h0EA7: data <= 32'hA5F25178;	13'h0EA8: data <= 32'hA60196D7;	13'h0EA9: data <= 32'hA610DC36;	13'h0EAA: data <= 32'hA6202194;	13'h0EAB: data <= 32'hA62F66F3;	13'h0EAC: data <= 32'hA63EAC52;	13'h0EAD: data <= 32'hA64DF1B1;	13'h0EAE: data <= 32'hA65D1FC5;	13'h0EAF: data <= 32'hA66C2E3B;	13'h0EB0: data <= 32'hA67B3CB2;	13'h0EB1: data <= 32'hA68A4B29;	13'h0EB2: data <= 32'hA699599F;	13'h0EB3: data <= 32'hA6A86816;	13'h0EB4: data <= 32'hA6B7768D;	13'h0EB5: data <= 32'hA6C68503;	13'h0EB6: data <= 32'hA6D5937A;	13'h0EB7: data <= 32'hA6E4A1F1;	13'h0EB8: data <= 32'hA6F3B067;	13'h0EB9: data <= 32'hA702BEDE;	13'h0EBA: data <= 32'hA711CD55;	13'h0EBB: data <= 32'hA720DBCB;	13'h0EBC: data <= 32'hA72FEA42;	13'h0EBD: data <= 32'hA73EF8B9;	13'h0EBE: data <= 32'hA74E072F;	13'h0EBF: data <= 32'hA75D15A6;	13'h0EC0: data <= 32'hA76C241D;	13'h0EC1: data <= 32'hA77B3293;	13'h0EC2: data <= 32'hA78A410A;	13'h0EC3: data <= 32'hA7994F81;	13'h0EC4: data <= 32'hA7A85DF7;	13'h0EC5: data <= 32'hA7B76C6E;	13'h0EC6: data <= 32'hA7C67AE5;	13'h0EC7: data <= 32'hA7D5895B;	13'h0EC8: data <= 32'hA7E497D2;	13'h0EC9: data <= 32'hA7F3A649;	13'h0ECA: data <= 32'hA802B4BF;	13'h0ECB: data <= 32'hA811C336;	13'h0ECC: data <= 32'hA820A9BE;	13'h0ECD: data <= 32'hA82E6EC4;	13'h0ECE: data <= 32'hA83C33C9;	13'h0ECF: data <= 32'hA849F8CF;	13'h0ED0: data <= 32'hA857BDD5;	13'h0ED1: data <= 32'hA86582DB;	13'h0ED2: data <= 32'hA87347E0;	13'h0ED3: data <= 32'hA8810CE6;	13'h0ED4: data <= 32'hA88ED1EC;	13'h0ED5: data <= 32'hA89C96F2;	13'h0ED6: data <= 32'hA8AA5BF7;	13'h0ED7: data <= 32'hA8B820FD;	13'h0ED8: data <= 32'hA8C5E603;	13'h0ED9: data <= 32'hA8D3AB08;	13'h0EDA: data <= 32'hA8E1700E;	13'h0EDB: data <= 32'hA8EF3514;	13'h0EDC: data <= 32'hA8FCFA1A;	13'h0EDD: data <= 32'hA90ABF1F;	13'h0EDE: data <= 32'hA9188425;	13'h0EDF: data <= 32'hA926492B;	13'h0EE0: data <= 32'hA9340E30;	13'h0EE1: data <= 32'hA941D336;	13'h0EE2: data <= 32'hA94F983C;	13'h0EE3: data <= 32'hA95D5D42;	13'h0EE4: data <= 32'hA96B2247;	13'h0EE5: data <= 32'hA978E74D;	13'h0EE6: data <= 32'hA986AC53;	13'h0EE7: data <= 32'hA9947159;	13'h0EE8: data <= 32'hA9A2365E;	13'h0EE9: data <= 32'hA9AFFB64;	13'h0EEA: data <= 32'hA9BDC06A;	13'h0EEB: data <= 32'hA9C9F59D;	13'h0EEC: data <= 32'hA9D5D1F7;	13'h0EED: data <= 32'hA9E1AE51;	13'h0EEE: data <= 32'hA9ED8AAB;	13'h0EEF: data <= 32'hA9F96704;	13'h0EF0: data <= 32'hAA05435E;	13'h0EF1: data <= 32'hAA111FB8;	13'h0EF2: data <= 32'hAA1CFC12;	13'h0EF3: data <= 32'hAA28D86C;	13'h0EF4: data <= 32'hAA34B4C6;	13'h0EF5: data <= 32'hAA409120;	13'h0EF6: data <= 32'hAA4C6D79;	13'h0EF7: data <= 32'hAA5849D3;	13'h0EF8: data <= 32'hAA64262D;	13'h0EF9: data <= 32'hAA700287;	13'h0EFA: data <= 32'hAA7BDEE1;	13'h0EFB: data <= 32'hAA87BB3B;	13'h0EFC: data <= 32'hAA939795;	13'h0EFD: data <= 32'hAA9F73EE;	13'h0EFE: data <= 32'hAAAB5048;	13'h0EFF: data <= 32'hAAB72CA2;	13'h0F00: data <= 32'hAAC308FC;	13'h0F01: data <= 32'hAACEE556;	13'h0F02: data <= 32'hAADAC1B0;	13'h0F03: data <= 32'hAAE69E0A;	13'h0F04: data <= 32'hAAF27A63;	13'h0F05: data <= 32'hAAFE56BD;	13'h0F06: data <= 32'hAB0A3317;	13'h0F07: data <= 32'hAB160F71;	13'h0F08: data <= 32'hAB21EBCB;	13'h0F09: data <= 32'hAB2C74B8;	13'h0F0A: data <= 32'hAB35BE30;	13'h0F0B: data <= 32'hAB3F07A8;	13'h0F0C: data <= 32'hAB485120;	13'h0F0D: data <= 32'hAB519A98;	13'h0F0E: data <= 32'hAB5AE40F;	13'h0F0F: data <= 32'hAB642D87;	13'h0F10: data <= 32'hAB6D76FF;	13'h0F11: data <= 32'hAB76C077;	13'h0F12: data <= 32'hAB8009EF;	13'h0F13: data <= 32'hAB895367;	13'h0F14: data <= 32'hAB929CDF;	13'h0F15: data <= 32'hAB9BE657;	13'h0F16: data <= 32'hABA52FCE;	13'h0F17: data <= 32'hABAE7946;	13'h0F18: data <= 32'hABB7C2BE;	13'h0F19: data <= 32'hABC10C36;	13'h0F1A: data <= 32'hABCA55AE;	13'h0F1B: data <= 32'hABD39F26;	13'h0F1C: data <= 32'hABDCE89E;	13'h0F1D: data <= 32'hABE63216;	13'h0F1E: data <= 32'hABEF7B8D;	13'h0F1F: data <= 32'hABF8C505;	13'h0F20: data <= 32'hAC020E7D;	13'h0F21: data <= 32'hAC0B57F5;	13'h0F22: data <= 32'hAC14A16D;	13'h0F23: data <= 32'hAC1DEAE5;	13'h0F24: data <= 32'hAC27345D;	13'h0F25: data <= 32'hAC307DD4;	13'h0F26: data <= 32'hAC39C74C;	13'h0F27: data <= 32'hAC42725E;	13'h0F28: data <= 32'hAC48D11A;	13'h0F29: data <= 32'hAC4F2FD6;	13'h0F2A: data <= 32'hAC558E92;	13'h0F2B: data <= 32'hAC5BED4F;	13'h0F2C: data <= 32'hAC624C0B;	13'h0F2D: data <= 32'hAC68AAC7;	13'h0F2E: data <= 32'hAC6F0983;	13'h0F2F: data <= 32'hAC75683F;	13'h0F30: data <= 32'hAC7BC6FB;	13'h0F31: data <= 32'hAC8225B7;	13'h0F32: data <= 32'hAC888473;	13'h0F33: data <= 32'hAC8EE32F;	13'h0F34: data <= 32'hAC9541EB;	13'h0F35: data <= 32'hAC9BA0A7;	13'h0F36: data <= 32'hACA1FF63;	13'h0F37: data <= 32'hACA85E1F;	13'h0F38: data <= 32'hACAEBCDB;	13'h0F39: data <= 32'hACB51B97;	13'h0F3A: data <= 32'hACBB7A53;	13'h0F3B: data <= 32'hACC1D90F;	13'h0F3C: data <= 32'hACC837CB;	13'h0F3D: data <= 32'hACCE9687;	13'h0F3E: data <= 32'hACD4F544;	13'h0F3F: data <= 32'hACDB5400;	13'h0F40: data <= 32'hACE1B2BC;	13'h0F41: data <= 32'hACE81178;	13'h0F42: data <= 32'hACEE7034;	13'h0F43: data <= 32'hACF4CEF0;	13'h0F44: data <= 32'hACFB2DAC;	13'h0F45: data <= 32'hAD018C68;	13'h0F46: data <= 32'hAD05EE01;	13'h0F47: data <= 32'hAD0A1CB0;	13'h0F48: data <= 32'hAD0E4B5F;	13'h0F49: data <= 32'hAD127A0F;	13'h0F4A: data <= 32'hAD16A8BE;	13'h0F4B: data <= 32'hAD1AD76D;	13'h0F4C: data <= 32'hAD1F061C;	13'h0F4D: data <= 32'hAD2334CB;	13'h0F4E: data <= 32'hAD27637B;	13'h0F4F: data <= 32'hAD2B922A;	13'h0F50: data <= 32'hAD2FC0D9;	13'h0F51: data <= 32'hAD33EF88;	13'h0F52: data <= 32'hAD381E37;	13'h0F53: data <= 32'hAD3C4CE6;	13'h0F54: data <= 32'hAD407B96;	13'h0F55: data <= 32'hAD44AA45;	13'h0F56: data <= 32'hAD48D8F4;	13'h0F57: data <= 32'hAD4D07A3;	13'h0F58: data <= 32'hAD513652;	13'h0F59: data <= 32'hAD556502;	13'h0F5A: data <= 32'hAD5993B1;	13'h0F5B: data <= 32'hAD5DC260;	13'h0F5C: data <= 32'hAD61F10F;	13'h0F5D: data <= 32'hAD661FBE;	13'h0F5E: data <= 32'hAD6A4E6E;	13'h0F5F: data <= 32'hAD6E7D1D;	13'h0F60: data <= 32'hAD72ABCC;	13'h0F61: data <= 32'hAD76DA7B;	13'h0F62: data <= 32'hAD7B092A;	13'h0F63: data <= 32'hAD7F37DA;	13'h0F64: data <= 32'hAD830CB0;	13'h0F65: data <= 32'hAD86A71F;	13'h0F66: data <= 32'hAD8A418F;	13'h0F67: data <= 32'hAD8DDBFE;	13'h0F68: data <= 32'hAD91766E;	13'h0F69: data <= 32'hAD9510DE;	13'h0F6A: data <= 32'hAD98AB4D;	13'h0F6B: data <= 32'hAD9C45BD;	13'h0F6C: data <= 32'hAD9FE02C;	13'h0F6D: data <= 32'hADA37A9C;	13'h0F6E: data <= 32'hADA7150B;	13'h0F6F: data <= 32'hADAAAF7B;	13'h0F70: data <= 32'hADAE49EA;	13'h0F71: data <= 32'hADB1E45A;	13'h0F72: data <= 32'hADB57EC9;	13'h0F73: data <= 32'hADB91939;	13'h0F74: data <= 32'hADBCB3A9;	13'h0F75: data <= 32'hADC04E18;	13'h0F76: data <= 32'hADC3E888;	13'h0F77: data <= 32'hADC782F7;	13'h0F78: data <= 32'hADCB1D67;	13'h0F79: data <= 32'hADCEB7D6;	13'h0F7A: data <= 32'hADD25246;	13'h0F7B: data <= 32'hADD5ECB5;	13'h0F7C: data <= 32'hADD98725;	13'h0F7D: data <= 32'hADDD2194;	13'h0F7E: data <= 32'hADE0BC04;	13'h0F7F: data <= 32'hADE45674;	13'h0F80: data <= 32'hADE7F0E3;	13'h0F81: data <= 32'hADEB8B53;	13'h0F82: data <= 32'hADEF7C47;	13'h0F83: data <= 32'hADF4343B;	13'h0F84: data <= 32'hADF8EC2E;	13'h0F85: data <= 32'hADFDA422;	13'h0F86: data <= 32'hAE025C16;	13'h0F87: data <= 32'hAE071409;	13'h0F88: data <= 32'hAE0BCBFD;	13'h0F89: data <= 32'hAE1083F1;	13'h0F8A: data <= 32'hAE153BE4;	13'h0F8B: data <= 32'hAE19F3D8;	13'h0F8C: data <= 32'hAE1EABCB;	13'h0F8D: data <= 32'hAE2363BF;	13'h0F8E: data <= 32'hAE281BB3;	13'h0F8F: data <= 32'hAE2CD3A6;	13'h0F90: data <= 32'hAE318B9A;	13'h0F91: data <= 32'hAE36438D;	13'h0F92: data <= 32'hAE3AFB81;	13'h0F93: data <= 32'hAE3FB375;	13'h0F94: data <= 32'hAE446B68;	13'h0F95: data <= 32'hAE49235C;	13'h0F96: data <= 32'hAE4DDB4F;	13'h0F97: data <= 32'hAE529343;	13'h0F98: data <= 32'hAE574B37;	13'h0F99: data <= 32'hAE5C032A;	13'h0F9A: data <= 32'hAE60BB1E;	13'h0F9B: data <= 32'hAE657311;	13'h0F9C: data <= 32'hAE6A2B05;	13'h0F9D: data <= 32'hAE6EE2F9;	13'h0F9E: data <= 32'hAE739AEC;	13'h0F9F: data <= 32'hAE7852E0;	13'h0FA0: data <= 32'hAE7D0AD3;	13'h0FA1: data <= 32'hAE84711D;	13'h0FA2: data <= 32'hAE8BD767;	13'h0FA3: data <= 32'hAE933DB0;	13'h0FA4: data <= 32'hAE9AA3FA;	13'h0FA5: data <= 32'hAEA20A44;	13'h0FA6: data <= 32'hAEA9708D;	13'h0FA7: data <= 32'hAEB0D6D7;	13'h0FA8: data <= 32'hAEB83D21;	13'h0FA9: data <= 32'hAEBFA36A;	13'h0FAA: data <= 32'hAEC709B4;	13'h0FAB: data <= 32'hAECE6FFE;	13'h0FAC: data <= 32'hAED5D647;	13'h0FAD: data <= 32'hAEDD3C91;	13'h0FAE: data <= 32'hAEE4A2DA;	13'h0FAF: data <= 32'hAEEC0924;	13'h0FB0: data <= 32'hAEF36F6E;	13'h0FB1: data <= 32'hAEFAD5B7;	13'h0FB2: data <= 32'hAF023C01;	13'h0FB3: data <= 32'hAF09A24B;	13'h0FB4: data <= 32'hAF110894;	13'h0FB5: data <= 32'hAF186EDE;	13'h0FB6: data <= 32'hAF1FD528;	13'h0FB7: data <= 32'hAF273B71;	13'h0FB8: data <= 32'hAF2EA1BB;	13'h0FB9: data <= 32'hAF360804;	13'h0FBA: data <= 32'hAF3D6E4E;	13'h0FBB: data <= 32'hAF44D498;	13'h0FBC: data <= 32'hAF4C3AE1;	13'h0FBD: data <= 32'hAF53A12B;	13'h0FBE: data <= 32'hAF5B0775;	13'h0FBF: data <= 32'hAF6531B6;	13'h0FC0: data <= 32'hAF708FC6;	13'h0FC1: data <= 32'hAF7BEDD7;	13'h0FC2: data <= 32'hAF874BE8;	13'h0FC3: data <= 32'hAF92A9F8;	13'h0FC4: data <= 32'hAF9E0809;	13'h0FC5: data <= 32'hAFA9661A;	13'h0FC6: data <= 32'hAFB4C42A;	13'h0FC7: data <= 32'hAFC0223B;	13'h0FC8: data <= 32'hAFCB804C;	13'h0FC9: data <= 32'hAFD6DE5D;	13'h0FCA: data <= 32'hAFE23C6D;	13'h0FCB: data <= 32'hAFED9A7E;	13'h0FCC: data <= 32'hAFF8F88F;	13'h0FCD: data <= 32'hB004569F;	13'h0FCE: data <= 32'hB00FB4B0;	13'h0FCF: data <= 32'hB01B12C1;	13'h0FD0: data <= 32'hB02670D1;	13'h0FD1: data <= 32'hB031CEE2;	13'h0FD2: data <= 32'hB03D2CF3;	13'h0FD3: data <= 32'hB0488B03;	13'h0FD4: data <= 32'hB053E914;	13'h0FD5: data <= 32'hB05F4725;	13'h0FD6: data <= 32'hB06AA535;	13'h0FD7: data <= 32'hB0760346;	13'h0FD8: data <= 32'hB0816157;	13'h0FD9: data <= 32'hB08CBF67;	13'h0FDA: data <= 32'hB0981D78;	13'h0FDB: data <= 32'hB0A37B89;	13'h0FDC: data <= 32'hB0AED999;	13'h0FDD: data <= 32'hB0BC22AA;	13'h0FDE: data <= 32'hB0CC5F1E;	13'h0FDF: data <= 32'hB0DC9B92;	13'h0FE0: data <= 32'hB0ECD805;	13'h0FE1: data <= 32'hB0FD1479;	13'h0FE2: data <= 32'hB10D50EC;	13'h0FE3: data <= 32'hB11D8D60;	13'h0FE4: data <= 32'hB12DC9D4;	13'h0FE5: data <= 32'hB13E0647;	13'h0FE6: data <= 32'hB14E42BB;	13'h0FE7: data <= 32'hB15E7F2E;	13'h0FE8: data <= 32'hB16EBBA2;	13'h0FE9: data <= 32'hB17EF816;	13'h0FEA: data <= 32'hB18F3489;	13'h0FEB: data <= 32'hB19F70FD;	13'h0FEC: data <= 32'hB1AFAD70;	13'h0FED: data <= 32'hB1BFE9E4;	13'h0FEE: data <= 32'hB1D02658;	13'h0FEF: data <= 32'hB1E062CB;	13'h0FF0: data <= 32'hB1F09F3F;	13'h0FF1: data <= 32'hB200DBB2;	13'h0FF2: data <= 32'hB2111826;	13'h0FF3: data <= 32'hB221549A;	13'h0FF4: data <= 32'hB231910D;	13'h0FF5: data <= 32'hB241CD81;	13'h0FF6: data <= 32'hB25209F4;	13'h0FF7: data <= 32'hB2624668;	13'h0FF8: data <= 32'hB27282DC;	13'h0FF9: data <= 32'hB282BF4F;	13'h0FFA: data <= 32'hB292FBC3;	13'h0FFB: data <= 32'hB2A3A607;	13'h0FFC: data <= 32'hB2B89A6E;	13'h0FFD: data <= 32'hB2CD8ED5;	13'h0FFE: data <= 32'hB2E2833C;	13'h0FFF: data <= 32'hB2F777A4;	13'h1000: data <= 32'hB30C6C0B;	13'h1001: data <= 32'hB3216072;	13'h1002: data <= 32'hB33654D9;	13'h1003: data <= 32'hB34B4940;	13'h1004: data <= 32'hB3603DA7;	13'h1005: data <= 32'hB375320F;	13'h1006: data <= 32'hB38A2676;	13'h1007: data <= 32'hB39F1ADD;	13'h1008: data <= 32'hB3B40F44;	13'h1009: data <= 32'hB3C903AB;	13'h100A: data <= 32'hB3DDF812;	13'h100B: data <= 32'hB3F2EC7A;	13'h100C: data <= 32'hB407E0E1;	13'h100D: data <= 32'hB41CD548;	13'h100E: data <= 32'hB431C9AF;	13'h100F: data <= 32'hB446BE16;	13'h1010: data <= 32'hB45BB27E;	13'h1011: data <= 32'hB470A6E5;	13'h1012: data <= 32'hB4859B4C;	13'h1013: data <= 32'hB49A8FB3;	13'h1014: data <= 32'hB4AF841A;	13'h1015: data <= 32'hB4C47881;	13'h1016: data <= 32'hB4D96CE9;	13'h1017: data <= 32'hB4EE6150;	13'h1018: data <= 32'hB50355B7;	13'h1019: data <= 32'hB5184A1E;	13'h101A: data <= 32'hB53051DA;	13'h101B: data <= 32'hB5492D90;	13'h101C: data <= 32'hB5620945;	13'h101D: data <= 32'hB57AE4FA;	13'h101E: data <= 32'hB593C0B0;	13'h101F: data <= 32'hB5AC9C65;	13'h1020: data <= 32'hB5C5781B;	13'h1021: data <= 32'hB5DE53D0;	13'h1022: data <= 32'hB5F72F85;	13'h1023: data <= 32'hB6100B3B;	13'h1024: data <= 32'hB628E6F0;	13'h1025: data <= 32'hB641C2A5;	13'h1026: data <= 32'hB65A9E5B;	13'h1027: data <= 32'hB6737A10;	13'h1028: data <= 32'hB68C55C6;	13'h1029: data <= 32'hB6A5317B;	13'h102A: data <= 32'hB6BE0D30;	13'h102B: data <= 32'hB6D6E8E6;	13'h102C: data <= 32'hB6EFC49B;	13'h102D: data <= 32'hB708A051;	13'h102E: data <= 32'hB7217C06;	13'h102F: data <= 32'hB73A57BB;	13'h1030: data <= 32'hB7533371;	13'h1031: data <= 32'hB76C0F26;	13'h1032: data <= 32'hB784EADB;	13'h1033: data <= 32'hB79DC691;	13'h1034: data <= 32'hB7B6A246;	13'h1035: data <= 32'hB7CF7DFC;	13'h1036: data <= 32'hB7E859B1;	13'h1037: data <= 32'hB8013566;	13'h1038: data <= 32'hB81BA06E;	13'h1039: data <= 32'hB837B3BE;	13'h103A: data <= 32'hB853C70E;	13'h103B: data <= 32'hB86FDA5E;	13'h103C: data <= 32'hB88BEDAE;	13'h103D: data <= 32'hB8A800FD;	13'h103E: data <= 32'hB8C4144D;	13'h103F: data <= 32'hB8E0279D;	13'h1040: data <= 32'hB8FC3AED;	13'h1041: data <= 32'hB9184E3C;	13'h1042: data <= 32'hB934618C;	13'h1043: data <= 32'hB95074DC;	13'h1044: data <= 32'hB96C882C;	13'h1045: data <= 32'hB9889B7C;	13'h1046: data <= 32'hB9A4AECB;	13'h1047: data <= 32'hB9C0C21B;	13'h1048: data <= 32'hB9DCD56B;	13'h1049: data <= 32'hB9F8E8BB;	13'h104A: data <= 32'hBA14FC0B;	13'h104B: data <= 32'hBA310F5A;	13'h104C: data <= 32'hBA4D22AA;	13'h104D: data <= 32'hBA6935FA;	13'h104E: data <= 32'hBA85494A;	13'h104F: data <= 32'hBAA15C9A;	13'h1050: data <= 32'hBABD6FE9;	13'h1051: data <= 32'hBAD98339;	13'h1052: data <= 32'hBAF59689;	13'h1053: data <= 32'hBB11A9D9;	13'h1054: data <= 32'hBB2DBD29;	13'h1055: data <= 32'hBB49D078;	13'h1056: data <= 32'hBB666291;	13'h1057: data <= 32'hBB852F32;	13'h1058: data <= 32'hBBA3FBD3;	13'h1059: data <= 32'hBBC2C875;	13'h105A: data <= 32'hBBE19516;	13'h105B: data <= 32'hBC0061B7;	13'h105C: data <= 32'hBC1F2E58;	13'h105D: data <= 32'hBC3DFAF9;	13'h105E: data <= 32'hBC5CC79A;	13'h105F: data <= 32'hBC7B943B;	13'h1060: data <= 32'hBC9A60DC;	13'h1061: data <= 32'hBCB92D7E;	13'h1062: data <= 32'hBCD7FA1F;	13'h1063: data <= 32'hBCF6C6C0;	13'h1064: data <= 32'hBD159361;	13'h1065: data <= 32'hBD346002;	13'h1066: data <= 32'hBD532CA3;	13'h1067: data <= 32'hBD71F944;	13'h1068: data <= 32'hBD90C5E5;	13'h1069: data <= 32'hBDAF9287;	13'h106A: data <= 32'hBDCE5F28;	13'h106B: data <= 32'hBDED2BC9;	13'h106C: data <= 32'hBE0BF86A;	13'h106D: data <= 32'hBE2AC50B;	13'h106E: data <= 32'hBE4991AC;	13'h106F: data <= 32'hBE685E4D;	13'h1070: data <= 32'hBE872AEF;	13'h1071: data <= 32'hBEA5F790;	13'h1072: data <= 32'hBEC4C431;	13'h1073: data <= 32'hBEE390D2;	13'h1074: data <= 32'hBF025D73;	13'h1075: data <= 32'hBF22AC17;	13'h1076: data <= 32'hBF432FFA;	13'h1077: data <= 32'hBF63B3DC;	13'h1078: data <= 32'hBF8437BE;	13'h1079: data <= 32'hBFA4BBA1;	13'h107A: data <= 32'hBFC53F83;	13'h107B: data <= 32'hBFE5C366;	13'h107C: data <= 32'hC0064748;	13'h107D: data <= 32'hC026CB2B;	13'h107E: data <= 32'hC0474F0D;	13'h107F: data <= 32'hC067D2EF;	13'h1080: data <= 32'hC08856D2;	13'h1081: data <= 32'hC0A8DAB4;	13'h1082: data <= 32'hC0C95E97;	13'h1083: data <= 32'hC0E9E279;	13'h1084: data <= 32'hC10A665B;	13'h1085: data <= 32'hC12AEA3E;	13'h1086: data <= 32'hC14B6E20;	13'h1087: data <= 32'hC16BF203;	13'h1088: data <= 32'hC18C75E5;	13'h1089: data <= 32'hC1ACF9C7;	13'h108A: data <= 32'hC1CD7DAA;	13'h108B: data <= 32'hC1EE018C;	13'h108C: data <= 32'hC20E856F;	13'h108D: data <= 32'hC22F0951;	13'h108E: data <= 32'hC24F8D34;	13'h108F: data <= 32'hC2701116;	13'h1090: data <= 32'hC29094F8;	13'h1091: data <= 32'hC2B118DB;	13'h1092: data <= 32'hC2D19CBD;	13'h1093: data <= 32'hC2F2500B;	13'h1094: data <= 32'hC313264A;	13'h1095: data <= 32'hC333FC88;	13'h1096: data <= 32'hC354D2C7;	13'h1097: data <= 32'hC375A906;	13'h1098: data <= 32'hC3967F44;	13'h1099: data <= 32'hC3B75583;	13'h109A: data <= 32'hC3D82BC1;	13'h109B: data <= 32'hC3F90200;	13'h109C: data <= 32'hC419D83F;	13'h109D: data <= 32'hC43AAE7D;	13'h109E: data <= 32'hC45B84BC;	13'h109F: data <= 32'hC47C5AFB;	13'h10A0: data <= 32'hC49D3139;	13'h10A1: data <= 32'hC4BE0778;	13'h10A2: data <= 32'hC4DEDDB7;	13'h10A3: data <= 32'hC4FFB3F5;	13'h10A4: data <= 32'hC5208A34;	13'h10A5: data <= 32'hC5416073;	13'h10A6: data <= 32'hC56236B1;	13'h10A7: data <= 32'hC5830CF0;	13'h10A8: data <= 32'hC5A3E32E;	13'h10A9: data <= 32'hC5C4B96D;	13'h10AA: data <= 32'hC5E58FAC;	13'h10AB: data <= 32'hC60665EA;	13'h10AC: data <= 32'hC6273C29;	13'h10AD: data <= 32'hC6481268;	13'h10AE: data <= 32'hC668E8A6;	13'h10AF: data <= 32'hC689BEE5;	13'h10B0: data <= 32'hC6AA9524;	13'h10B1: data <= 32'hC6CB2C7E;	13'h10B2: data <= 32'hC6EB1C20;	13'h10B3: data <= 32'hC70B0BC3;	13'h10B4: data <= 32'hC72AFB66;	13'h10B5: data <= 32'hC74AEB09;	13'h10B6: data <= 32'hC76ADAAB;	13'h10B7: data <= 32'hC78ACA4E;	13'h10B8: data <= 32'hC7AAB9F1;	13'h10B9: data <= 32'hC7CAA994;	13'h10BA: data <= 32'hC7EA9936;	13'h10BB: data <= 32'hC80A88D9;	13'h10BC: data <= 32'hC82A787C;	13'h10BD: data <= 32'hC84A681F;	13'h10BE: data <= 32'hC86A57C1;	13'h10BF: data <= 32'hC88A4764;	13'h10C0: data <= 32'hC8AA3707;	13'h10C1: data <= 32'hC8CA26AA;	13'h10C2: data <= 32'hC8EA164C;	13'h10C3: data <= 32'hC90A05EF;	13'h10C4: data <= 32'hC929F592;	13'h10C5: data <= 32'hC949E535;	13'h10C6: data <= 32'hC969D4D8;	13'h10C7: data <= 32'hC989C47A;	13'h10C8: data <= 32'hC9A9B41D;	13'h10C9: data <= 32'hC9C9A3C0;	13'h10CA: data <= 32'hC9E99363;	13'h10CB: data <= 32'hCA098305;	13'h10CC: data <= 32'hCA2972A8;	13'h10CD: data <= 32'hCA49624B;	13'h10CE: data <= 32'hCA6951EE;	13'h10CF: data <= 32'hCA894190;	13'h10D0: data <= 32'hCAA7F711;	13'h10D1: data <= 32'hCAC6A2C0;	13'h10D2: data <= 32'hCAE54E70;	13'h10D3: data <= 32'hCB03FA1F;	13'h10D4: data <= 32'hCB22A5CF;	13'h10D5: data <= 32'hCB41517E;	13'h10D6: data <= 32'hCB5FFD2D;	13'h10D7: data <= 32'hCB7EA8DD;	13'h10D8: data <= 32'hCB9D548C;	13'h10D9: data <= 32'hCBBC003C;	13'h10DA: data <= 32'hCBDAABEB;	13'h10DB: data <= 32'hCBF9579A;	13'h10DC: data <= 32'hCC18034A;	13'h10DD: data <= 32'hCC36AEF9;	13'h10DE: data <= 32'hCC555AA9;	13'h10DF: data <= 32'hCC740658;	13'h10E0: data <= 32'hCC92B208;	13'h10E1: data <= 32'hCCB15DB7;	13'h10E2: data <= 32'hCCD00966;	13'h10E3: data <= 32'hCCEEB516;	13'h10E4: data <= 32'hCD0D60C5;	13'h10E5: data <= 32'hCD2C0C75;	13'h10E6: data <= 32'hCD4AB824;	13'h10E7: data <= 32'hCD6963D4;	13'h10E8: data <= 32'hCD880F83;	13'h10E9: data <= 32'hCDA6BB32;	13'h10EA: data <= 32'hCDC566E2;	13'h10EB: data <= 32'hCDE41291;	13'h10EC: data <= 32'hCE02BE41;	13'h10ED: data <= 32'hCE2169F0;	13'h10EE: data <= 32'hCE3F4C4C;	13'h10EF: data <= 32'hCE5CC9FF;	13'h10F0: data <= 32'hCE7A47B1;	13'h10F1: data <= 32'hCE97C564;	13'h10F2: data <= 32'hCEB54316;	13'h10F3: data <= 32'hCED2C0C9;	13'h10F4: data <= 32'hCEF03E7B;	13'h10F5: data <= 32'hCF0DBC2E;	13'h10F6: data <= 32'hCF2B39E0;	13'h10F7: data <= 32'hCF48B793;	13'h10F8: data <= 32'hCF663545;	13'h10F9: data <= 32'hCF83B2F8;	13'h10FA: data <= 32'hCFA130AA;	13'h10FB: data <= 32'hCFBEAE5D;	13'h10FC: data <= 32'hCFDC2C0F;	13'h10FD: data <= 32'hCFF9A9C2;	13'h10FE: data <= 32'hD0172774;	13'h10FF: data <= 32'hD034A527;	13'h1100: data <= 32'hD05222D9;	13'h1101: data <= 32'hD06FA08C;	13'h1102: data <= 32'hD08D1E3F;	13'h1103: data <= 32'hD0AA9BF1;	13'h1104: data <= 32'hD0C819A4;	13'h1105: data <= 32'hD0E59756;	13'h1106: data <= 32'hD1031509;	13'h1107: data <= 32'hD12092BB;	13'h1108: data <= 32'hD13E106E;	13'h1109: data <= 32'hD15B8E20;	13'h110A: data <= 32'hD1790BD3;	13'h110B: data <= 32'hD1968985;	13'h110C: data <= 32'hD1B39B66;	13'h110D: data <= 32'hD1CFF09A;	13'h110E: data <= 32'hD1EC45CD;	13'h110F: data <= 32'hD2089B00;	13'h1110: data <= 32'hD224F033;	13'h1111: data <= 32'hD2414567;	13'h1112: data <= 32'hD25D9A9A;	13'h1113: data <= 32'hD279EFCD;	13'h1114: data <= 32'hD2964500;	13'h1115: data <= 32'hD2B29A33;	13'h1116: data <= 32'hD2CEEF67;	13'h1117: data <= 32'hD2EB449A;	13'h1118: data <= 32'hD30799CD;	13'h1119: data <= 32'hD323EF00;	13'h111A: data <= 32'hD3404434;	13'h111B: data <= 32'hD35C9967;	13'h111C: data <= 32'hD378EE9A;	13'h111D: data <= 32'hD39543CD;	13'h111E: data <= 32'hD3B19900;	13'h111F: data <= 32'hD3CDEE34;	13'h1120: data <= 32'hD3EA4367;	13'h1121: data <= 32'hD406989A;	13'h1122: data <= 32'hD422EDCD;	13'h1123: data <= 32'hD43F4300;	13'h1124: data <= 32'hD45B9834;	13'h1125: data <= 32'hD477ED67;	13'h1126: data <= 32'hD494429A;	13'h1127: data <= 32'hD4B097CD;	13'h1128: data <= 32'hD4CCED01;	13'h1129: data <= 32'hD4E94234;	13'h112A: data <= 32'hD5058BC1;	13'h112B: data <= 32'hD52120C8;	13'h112C: data <= 32'hD53CB5CF;	13'h112D: data <= 32'hD5584AD5;	13'h112E: data <= 32'hD573DFDC;	13'h112F: data <= 32'hD58F74E2;	13'h1130: data <= 32'hD5AB09E9;	13'h1131: data <= 32'hD5C69EF0;	13'h1132: data <= 32'hD5E233F6;	13'h1133: data <= 32'hD5FDC8FD;	13'h1134: data <= 32'hD6195E04;	13'h1135: data <= 32'hD634F30A;	13'h1136: data <= 32'hD6508811;	13'h1137: data <= 32'hD66C1D17;	13'h1138: data <= 32'hD687B21E;	13'h1139: data <= 32'hD6A34725;	13'h113A: data <= 32'hD6BEDC2B;	13'h113B: data <= 32'hD6DA7132;	13'h113C: data <= 32'hD6F60639;	13'h113D: data <= 32'hD7119B3F;	13'h113E: data <= 32'hD72D3046;	13'h113F: data <= 32'hD748C54C;	13'h1140: data <= 32'hD7645A53;	13'h1141: data <= 32'hD77FEF5A;	13'h1142: data <= 32'hD79B8460;	13'h1143: data <= 32'hD7B71967;	13'h1144: data <= 32'hD7D2AE6D;	13'h1145: data <= 32'hD7EE4374;	13'h1146: data <= 32'hD809D87B;	13'h1147: data <= 32'hD8256D81;	13'h1148: data <= 32'hD8410288;	13'h1149: data <= 32'hD85D0C07;	13'h114A: data <= 32'hD8793ACB;	13'h114B: data <= 32'hD895698F;	13'h114C: data <= 32'hD8B19853;	13'h114D: data <= 32'hD8CDC716;	13'h114E: data <= 32'hD8E9F5DA;	13'h114F: data <= 32'hD906249E;	13'h1150: data <= 32'hD9225362;	13'h1151: data <= 32'hD93E8226;	13'h1152: data <= 32'hD95AB0EA;	13'h1153: data <= 32'hD976DFAE;	13'h1154: data <= 32'hD9930E72;	13'h1155: data <= 32'hD9AF3D36;	13'h1156: data <= 32'hD9CB6BFA;	13'h1157: data <= 32'hD9E79ABE;	13'h1158: data <= 32'hDA03C982;	13'h1159: data <= 32'hDA1FF846;	13'h115A: data <= 32'hDA3C270A;	13'h115B: data <= 32'hDA5855CE;	13'h115C: data <= 32'hDA748492;	13'h115D: data <= 32'hDA90B355;	13'h115E: data <= 32'hDAACE219;	13'h115F: data <= 32'hDAC910DD;	13'h1160: data <= 32'hDAE53FA1;	13'h1161: data <= 32'hDB016E65;	13'h1162: data <= 32'hDB1D9D29;	13'h1163: data <= 32'hDB39CBED;	13'h1164: data <= 32'hDB55FAB1;	13'h1165: data <= 32'hDB722975;	13'h1166: data <= 32'hDB8E5839;	13'h1167: data <= 32'hDBABD56C;	13'h1168: data <= 32'hDBCAE3F0;	13'h1169: data <= 32'hDBE9F275;	13'h116A: data <= 32'hDC0900F9;	13'h116B: data <= 32'hDC280F7E;	13'h116C: data <= 32'hDC471E02;	13'h116D: data <= 32'hDC662C87;	13'h116E: data <= 32'hDC853B0B;	13'h116F: data <= 32'hDCA44990;	13'h1170: data <= 32'hDCC35814;	13'h1171: data <= 32'hDCE26698;	13'h1172: data <= 32'hDD01751D;	13'h1173: data <= 32'hDD2083A1;	13'h1174: data <= 32'hDD3F9226;	13'h1175: data <= 32'hDD5EA0AA;	13'h1176: data <= 32'hDD7DAF2F;	13'h1177: data <= 32'hDD9CBDB3;	13'h1178: data <= 32'hDDBBCC38;	13'h1179: data <= 32'hDDDADABC;	13'h117A: data <= 32'hDDF9E941;	13'h117B: data <= 32'hDE18F7C5;	13'h117C: data <= 32'hDE38064A;	13'h117D: data <= 32'hDE5714CE;	13'h117E: data <= 32'hDE762353;	13'h117F: data <= 32'hDE9531D7;	13'h1180: data <= 32'hDEB4405C;	13'h1181: data <= 32'hDED34EE0;	13'h1182: data <= 32'hDEF25D65;	13'h1183: data <= 32'hDF116BE9;	13'h1184: data <= 32'hDF307A6E;	13'h1185: data <= 32'hDF505818;	13'h1186: data <= 32'hDF74BDCB;	13'h1187: data <= 32'hDF99237E;	13'h1188: data <= 32'hDFBD8931;	13'h1189: data <= 32'hDFE1EEE4;	13'h118A: data <= 32'hE0065497;	13'h118B: data <= 32'hE02ABA4A;	13'h118C: data <= 32'hE04F1FFD;	13'h118D: data <= 32'hE07385B0;	13'h118E: data <= 32'hE097EB63;	13'h118F: data <= 32'hE0BC5116;	13'h1190: data <= 32'hE0E0B6C9;	13'h1191: data <= 32'hE1051C7C;	13'h1192: data <= 32'hE129822F;	13'h1193: data <= 32'hE14DE7E2;	13'h1194: data <= 32'hE1724D95;	13'h1195: data <= 32'hE196B348;	13'h1196: data <= 32'hE1BB18FB;	13'h1197: data <= 32'hE1DF7EAE;	13'h1198: data <= 32'hE203E461;	13'h1199: data <= 32'hE2284A14;	13'h119A: data <= 32'hE24CAFC7;	13'h119B: data <= 32'hE271157A;	13'h119C: data <= 32'hE2957B2D;	13'h119D: data <= 32'hE2B9E0E0;	13'h119E: data <= 32'hE2DE4693;	13'h119F: data <= 32'hE302AC46;	13'h11A0: data <= 32'hE32711F9;	13'h11A1: data <= 32'hE34B77AC;	13'h11A2: data <= 32'hE36FDD5F;	13'h11A3: data <= 32'hE3944312;	13'h11A4: data <= 32'hE3BED417;	13'h11A5: data <= 32'hE3EA7F22;	13'h11A6: data <= 32'hE4162A2D;	13'h11A7: data <= 32'hE441D538;	13'h11A8: data <= 32'hE46D8043;	13'h11A9: data <= 32'hE4992B4E;	13'h11AA: data <= 32'hE4C4D659;	13'h11AB: data <= 32'hE4F08163;	13'h11AC: data <= 32'hE51C2C6E;	13'h11AD: data <= 32'hE547D779;	13'h11AE: data <= 32'hE5738284;	13'h11AF: data <= 32'hE59F2D8F;	13'h11B0: data <= 32'hE5CAD89A;	13'h11B1: data <= 32'hE5F683A5;	13'h11B2: data <= 32'hE6222EB0;	13'h11B3: data <= 32'hE64DD9BB;	13'h11B4: data <= 32'hE67984C6;	13'h11B5: data <= 32'hE6A52FD1;	13'h11B6: data <= 32'hE6D0DADB;	13'h11B7: data <= 32'hE6FC85E6;	13'h11B8: data <= 32'hE72830F1;	13'h11B9: data <= 32'hE753DBFC;	13'h11BA: data <= 32'hE77F8707;	13'h11BB: data <= 32'hE7AB3212;	13'h11BC: data <= 32'hE7D6DD1D;	13'h11BD: data <= 32'hE8028828;	13'h11BE: data <= 32'hE82E3333;	13'h11BF: data <= 32'hE859DE3E;	13'h11C0: data <= 32'hE8858949;	13'h11C1: data <= 32'hE8B13453;	13'h11C2: data <= 32'hE8E1BD42;	13'h11C3: data <= 32'hE916546D;	13'h11C4: data <= 32'hE94AEB98;	13'h11C5: data <= 32'hE97F82C4;	13'h11C6: data <= 32'hE9B419EF;	13'h11C7: data <= 32'hE9E8B11A;	13'h11C8: data <= 32'hEA1D4846;	13'h11C9: data <= 32'hEA51DF71;	13'h11CA: data <= 32'hEA86769C;	13'h11CB: data <= 32'hEABB0DC8;	13'h11CC: data <= 32'hEAEFA4F3;	13'h11CD: data <= 32'hEB243C1E;	13'h11CE: data <= 32'hEB58D34A;	13'h11CF: data <= 32'hEB8D6A75;	13'h11D0: data <= 32'hEBC201A0;	13'h11D1: data <= 32'hEBF698CC;	13'h11D2: data <= 32'hEC2B2FF7;	13'h11D3: data <= 32'hEC5FC722;	13'h11D4: data <= 32'hEC945E4E;	13'h11D5: data <= 32'hECC8F579;	13'h11D6: data <= 32'hECFD8CA4;	13'h11D7: data <= 32'hED3223D0;	13'h11D8: data <= 32'hED66BAFB;	13'h11D9: data <= 32'hED9B5227;	13'h11DA: data <= 32'hEDCFE952;	13'h11DB: data <= 32'hEE04807D;	13'h11DC: data <= 32'hEE3917A9;	13'h11DD: data <= 32'hEE6DAED4;	13'h11DE: data <= 32'hEEA245FF;	13'h11DF: data <= 32'hEED6DD2B;	13'h11E0: data <= 32'hEF0DE89B;	13'h11E1: data <= 32'hEF4C9F61;	13'h11E2: data <= 32'hEF8B5627;	13'h11E3: data <= 32'hEFCA0CED;	13'h11E4: data <= 32'hF008C3B3;	13'h11E5: data <= 32'hF0477A7A;	13'h11E6: data <= 32'hF0863140;	13'h11E7: data <= 32'hF0C4E806;	13'h11E8: data <= 32'hF1039ECC;	13'h11E9: data <= 32'hF1425593;	13'h11EA: data <= 32'hF1810C59;	13'h11EB: data <= 32'hF1BFC31F;	13'h11EC: data <= 32'hF1FE79E5;	13'h11ED: data <= 32'hF23D30AB;	13'h11EE: data <= 32'hF27BE772;	13'h11EF: data <= 32'hF2BA9E38;	13'h11F0: data <= 32'hF2F954FE;	13'h11F1: data <= 32'hF3380BC4;	13'h11F2: data <= 32'hF376C28B;	13'h11F3: data <= 32'hF3B57951;	13'h11F4: data <= 32'hF3F43017;	13'h11F5: data <= 32'hF432E6DD;	13'h11F6: data <= 32'hF4719DA3;	13'h11F7: data <= 32'hF4B0546A;	13'h11F8: data <= 32'hF4EF0B30;	13'h11F9: data <= 32'hF52DC1F6;	13'h11FA: data <= 32'hF56C78BC;	13'h11FB: data <= 32'hF5AB2F83;	13'h11FC: data <= 32'hF5E9E649;	13'h11FD: data <= 32'hF6289D0F;	13'h11FE: data <= 32'hF66753D5;	13'h11FF: data <= 32'hF6AFAC18;	13'h1200: data <= 32'hF6F8A36B;	13'h1201: data <= 32'hF7419ABE;	13'h1202: data <= 32'hF78A9211;	13'h1203: data <= 32'hF7D38964;	13'h1204: data <= 32'hF81C80B6;	13'h1205: data <= 32'hF8657809;	13'h1206: data <= 32'hF8AE6F5C;	13'h1207: data <= 32'hF8F766AF;	13'h1208: data <= 32'hF9405E02;	13'h1209: data <= 32'hF9895555;	13'h120A: data <= 32'hF9D24CA8;	13'h120B: data <= 32'hFA1B43FB;	13'h120C: data <= 32'hFA643B4E;	13'h120D: data <= 32'hFAAD32A1;	13'h120E: data <= 32'hFAF629F4;	13'h120F: data <= 32'hFB3F2146;	13'h1210: data <= 32'hFB881899;	13'h1211: data <= 32'hFBD10FEC;	13'h1212: data <= 32'hFC1A073F;	13'h1213: data <= 32'hFC62FE92;	13'h1214: data <= 32'hFCABF5E5;	13'h1215: data <= 32'hFCF4ED38;	13'h1216: data <= 32'hFD3DE48B;	13'h1217: data <= 32'hFD86DBDE;	13'h1218: data <= 32'hFDCFD331;	13'h1219: data <= 32'hFE18CA84;	13'h121A: data <= 32'hFE61C1D6;	13'h121B: data <= 32'hFEAAB929;	13'h121C: data <= 32'hFEF3B07C;	13'h121D: data <= 32'hFF426A4F;	13'h121E: data <= 32'hFF946EB4;	13'h121F: data <= 32'hFFE67319;	13'h1220: data <= 32'h0038777D;	13'h1221: data <= 32'h008A7BE2;	13'h1222: data <= 32'h00DC8047;	13'h1223: data <= 32'h012E84AC;	13'h1224: data <= 32'h01808910;	13'h1225: data <= 32'h01D28D75;	13'h1226: data <= 32'h022491DA;	13'h1227: data <= 32'h0276963F;	13'h1228: data <= 32'h02C89AA4;	13'h1229: data <= 32'h031A9F09;	13'h122A: data <= 32'h036CA36E;	13'h122B: data <= 32'h03BEA7D3;	13'h122C: data <= 32'h0410AC38;	13'h122D: data <= 32'h0462B09D;	13'h122E: data <= 32'h04B4B502;	13'h122F: data <= 32'h0506B967;	13'h1230: data <= 32'h0558BDCC;	13'h1231: data <= 32'h05AAC231;	13'h1232: data <= 32'h05FCC695;	13'h1233: data <= 32'h064ECAFA;	13'h1234: data <= 32'h06A0CF5F;	13'h1235: data <= 32'h06F2D3C4;	13'h1236: data <= 32'h0744D829;	13'h1237: data <= 32'h0796DC8E;	13'h1238: data <= 32'h07E8E0F3;	13'h1239: data <= 32'h083AE558;	13'h123A: data <= 32'h088CE9BD;	13'h123B: data <= 32'h08E16B0D;	13'h123C: data <= 32'h093AE635;	13'h123D: data <= 32'h0994615C;	13'h123E: data <= 32'h09EDDC84;	13'h123F: data <= 32'h0A4757AB;	13'h1240: data <= 32'h0AA0D2D3;	13'h1241: data <= 32'h0AFA4DFA;	13'h1242: data <= 32'h0B53C922;	13'h1243: data <= 32'h0BAD4449;	13'h1244: data <= 32'h0C06BF71;	13'h1245: data <= 32'h0C603A98;	13'h1246: data <= 32'h0CB9B5C0;	13'h1247: data <= 32'h0D1330E7;	13'h1248: data <= 32'h0D6CAC0F;	13'h1249: data <= 32'h0DC62736;	13'h124A: data <= 32'h0E1FA25E;	13'h124B: data <= 32'h0E791D85;	13'h124C: data <= 32'h0ED298AD;	13'h124D: data <= 32'h0F2C13D4;	13'h124E: data <= 32'h0F858EFC;	13'h124F: data <= 32'h0FDF0A23;	13'h1250: data <= 32'h1038854B;	13'h1251: data <= 32'h10920072;	13'h1252: data <= 32'h10EB7B9A;	13'h1253: data <= 32'h1144F6C1;	13'h1254: data <= 32'h119E71E9;	13'h1255: data <= 32'h11F7ED10;	13'h1256: data <= 32'h12516838;	13'h1257: data <= 32'h12AAE35F;	13'h1258: data <= 32'h13045E87;	13'h1259: data <= 32'h135E0148;	13'h125A: data <= 32'h13BC9738;	13'h125B: data <= 32'h141B2D28;	13'h125C: data <= 32'h1479C318;	13'h125D: data <= 32'h14D85909;	13'h125E: data <= 32'h1536EEF9;	13'h125F: data <= 32'h159584E9;	13'h1260: data <= 32'h15F41AD9;	13'h1261: data <= 32'h1652B0C9;	13'h1262: data <= 32'h16B146B9;	13'h1263: data <= 32'h170FDCA9;	13'h1264: data <= 32'h176E729A;	13'h1265: data <= 32'h17CD088A;	13'h1266: data <= 32'h182B9E7A;	13'h1267: data <= 32'h188A346A;	13'h1268: data <= 32'h18E8CA5A;	13'h1269: data <= 32'h1947604A;	13'h126A: data <= 32'h19A5F63A;	13'h126B: data <= 32'h1A048C2B;	13'h126C: data <= 32'h1A63221B;	13'h126D: data <= 32'h1AC1B80B;	13'h126E: data <= 32'h1B204DFB;	13'h126F: data <= 32'h1B7EE3EB;	13'h1270: data <= 32'h1BDD79DB;	13'h1271: data <= 32'h1C3C0FCB;	13'h1272: data <= 32'h1C9AA5BC;	13'h1273: data <= 32'h1CF93BAC;	13'h1274: data <= 32'h1D57D19C;	13'h1275: data <= 32'h1DB6678C;	13'h1276: data <= 32'h1E14FD7C;	13'h1277: data <= 32'h1E73936C;	13'h1278: data <= 32'h1ED398BD;	13'h1279: data <= 32'h1F3427D2;	13'h127A: data <= 32'h1F94B6E7;	13'h127B: data <= 32'h1FF545FC;	13'h127C: data <= 32'h2055D511;	13'h127D: data <= 32'h20B66425;	13'h127E: data <= 32'h2116F33A;	13'h127F: data <= 32'h2177824F;	13'h1280: data <= 32'h21D81164;	13'h1281: data <= 32'h2238A079;	13'h1282: data <= 32'h22992F8E;	13'h1283: data <= 32'h22F9BEA3;	13'h1284: data <= 32'h235A4DB8;	13'h1285: data <= 32'h23BADCCD;	13'h1286: data <= 32'h241B6BE1;	13'h1287: data <= 32'h247BFAF6;	13'h1288: data <= 32'h24DC8A0B;	13'h1289: data <= 32'h253D1920;	13'h128A: data <= 32'h259DA835;	13'h128B: data <= 32'h25FE374A;	13'h128C: data <= 32'h265EC65F;	13'h128D: data <= 32'h26BF5574;	13'h128E: data <= 32'h271FE489;	13'h128F: data <= 32'h2780739D;	13'h1290: data <= 32'h27E102B2;	13'h1291: data <= 32'h284191C7;	13'h1292: data <= 32'h28A220DC;	13'h1293: data <= 32'h2902AFF1;	13'h1294: data <= 32'h29633F06;	13'h1295: data <= 32'h29C3CE1B;	13'h1296: data <= 32'h2A23C5C7;	13'h1297: data <= 32'h2A82EFF6;	13'h1298: data <= 32'h2AE21A26;	13'h1299: data <= 32'h2B414456;	13'h129A: data <= 32'h2BA06E86;	13'h129B: data <= 32'h2BFF98B6;	13'h129C: data <= 32'h2C5EC2E6;	13'h129D: data <= 32'h2CBDED15;	13'h129E: data <= 32'h2D1D1745;	13'h129F: data <= 32'h2D7C4175;	13'h12A0: data <= 32'h2DDB6BA5;	13'h12A1: data <= 32'h2E3A95D5;	13'h12A2: data <= 32'h2E99C005;	13'h12A3: data <= 32'h2EF8EA34;	13'h12A4: data <= 32'h2F581464;	13'h12A5: data <= 32'h2FB73E94;	13'h12A6: data <= 32'h301668C4;	13'h12A7: data <= 32'h307592F4;	13'h12A8: data <= 32'h30D4BD24;	13'h12A9: data <= 32'h3133E753;	13'h12AA: data <= 32'h31931183;	13'h12AB: data <= 32'h31F23BB3;	13'h12AC: data <= 32'h325165E3;	13'h12AD: data <= 32'h32B09013;	13'h12AE: data <= 32'h330FBA43;	13'h12AF: data <= 32'h336EE472;	13'h12B0: data <= 32'h33CE0EA2;	13'h12B1: data <= 32'h342D38D2;	13'h12B2: data <= 32'h348C6302;	13'h12B3: data <= 32'h34EB8D32;	13'h12B4: data <= 32'h354A4792;	13'h12B5: data <= 32'h35A5D752;	13'h12B6: data <= 32'h36016713;	13'h12B7: data <= 32'h365CF6D3;	13'h12B8: data <= 32'h36B88693;	13'h12B9: data <= 32'h37141654;	13'h12BA: data <= 32'h376FA614;	13'h12BB: data <= 32'h37CB35D4;	13'h12BC: data <= 32'h3826C594;	13'h12BD: data <= 32'h38825555;	13'h12BE: data <= 32'h38DDE515;	13'h12BF: data <= 32'h393974D5;	13'h12C0: data <= 32'h39950495;	13'h12C1: data <= 32'h39F09456;	13'h12C2: data <= 32'h3A4C2416;	13'h12C3: data <= 32'h3AA7B3D6;	13'h12C4: data <= 32'h3B034397;	13'h12C5: data <= 32'h3B5ED357;	13'h12C6: data <= 32'h3BBA6317;	13'h12C7: data <= 32'h3C15F2D7;	13'h12C8: data <= 32'h3C718298;	13'h12C9: data <= 32'h3CCD1258;	13'h12CA: data <= 32'h3D28A218;	13'h12CB: data <= 32'h3D8431D9;	13'h12CC: data <= 32'h3DDFC199;	13'h12CD: data <= 32'h3E3B5159;	13'h12CE: data <= 32'h3E96E119;	13'h12CF: data <= 32'h3EF270DA;	13'h12D0: data <= 32'h3F4E009A;	13'h12D1: data <= 32'h3FA9905A;	13'h12D2: data <= 32'h4005201B;	13'h12D3: data <= 32'h405C2454;	13'h12D4: data <= 32'h40B225FE;	13'h12D5: data <= 32'h410827A7;	13'h12D6: data <= 32'h415E2951;	13'h12D7: data <= 32'h41B42AFA;	13'h12D8: data <= 32'h420A2CA4;	13'h12D9: data <= 32'h42602E4E;	13'h12DA: data <= 32'h42B62FF7;	13'h12DB: data <= 32'h430C31A1;	13'h12DC: data <= 32'h4362334A;	13'h12DD: data <= 32'h43B834F4;	13'h12DE: data <= 32'h440E369E;	13'h12DF: data <= 32'h44643847;	13'h12E0: data <= 32'h44BA39F1;	13'h12E1: data <= 32'h45103B9A;	13'h12E2: data <= 32'h45663D44;	13'h12E3: data <= 32'h45BC3EEE;	13'h12E4: data <= 32'h46124097;	13'h12E5: data <= 32'h46684241;	13'h12E6: data <= 32'h46BE43EA;	13'h12E7: data <= 32'h47144594;	13'h12E8: data <= 32'h476A473E;	13'h12E9: data <= 32'h47C048E7;	13'h12EA: data <= 32'h48164A91;	13'h12EB: data <= 32'h486C4C3B;	13'h12EC: data <= 32'h48C24DE4;	13'h12ED: data <= 32'h49184F8E;	13'h12EE: data <= 32'h496E5137;	13'h12EF: data <= 32'h49C452E1;	13'h12F0: data <= 32'h4A1A548B;	13'h12F1: data <= 32'h4A6C509E;	13'h12F2: data <= 32'h4ABA83AB;	13'h12F3: data <= 32'h4B08B6B8;	13'h12F4: data <= 32'h4B56E9C6;	13'h12F5: data <= 32'h4BA51CD3;	13'h12F6: data <= 32'h4BF34FE0;	13'h12F7: data <= 32'h4C4182EE;	13'h12F8: data <= 32'h4C8FB5FB;	13'h12F9: data <= 32'h4CDDE908;	13'h12FA: data <= 32'h4D2C1C15;	13'h12FB: data <= 32'h4D7A4F23;	13'h12FC: data <= 32'h4DC88230;	13'h12FD: data <= 32'h4E16B53D;	13'h12FE: data <= 32'h4E64E84B;	13'h12FF: data <= 32'h4EB31B58;	13'h1300: data <= 32'h4F014E65;	13'h1301: data <= 32'h4F4F8173;	13'h1302: data <= 32'h4F9DB480;	13'h1303: data <= 32'h4FEBE78D;	13'h1304: data <= 32'h503A1A9A;	13'h1305: data <= 32'h50884DA8;	13'h1306: data <= 32'h50D680B5;	13'h1307: data <= 32'h5124B3C2;	13'h1308: data <= 32'h5172E6D0;	13'h1309: data <= 32'h51C119DD;	13'h130A: data <= 32'h520F4CEA;	13'h130B: data <= 32'h525D7FF8;	13'h130C: data <= 32'h52ABB305;	13'h130D: data <= 32'h52F9E612;	13'h130E: data <= 32'h5348191F;	13'h130F: data <= 32'h5394642B;	13'h1310: data <= 32'h53D99A9F;	13'h1311: data <= 32'h541ED113;	13'h1312: data <= 32'h54640787;	13'h1313: data <= 32'h54A93DFB;	13'h1314: data <= 32'h54EE746F;	13'h1315: data <= 32'h5533AAE3;	13'h1316: data <= 32'h5578E157;	13'h1317: data <= 32'h55BE17CB;	13'h1318: data <= 32'h56034E3F;	13'h1319: data <= 32'h564884B3;	13'h131A: data <= 32'h568DBB27;	13'h131B: data <= 32'h56D2F19B;	13'h131C: data <= 32'h5718280F;	13'h131D: data <= 32'h575D5E83;	13'h131E: data <= 32'h57A294F7;	13'h131F: data <= 32'h57E7CB6B;	13'h1320: data <= 32'h582D01DF;	13'h1321: data <= 32'h58723853;	13'h1322: data <= 32'h58B76EC7;	13'h1323: data <= 32'h58FCA53B;	13'h1324: data <= 32'h5941DBAF;	13'h1325: data <= 32'h59871223;	13'h1326: data <= 32'h59CC4897;	13'h1327: data <= 32'h5A117F0B;	13'h1328: data <= 32'h5A56B57F;	13'h1329: data <= 32'h5A9BEBF3;	13'h132A: data <= 32'h5AE12267;	13'h132B: data <= 32'h5B2658DB;	13'h132C: data <= 32'h5B6B8F4F;	13'h132D: data <= 32'h5BB0C5C3;	13'h132E: data <= 32'h5BEDF8B1;	13'h132F: data <= 32'h5C2A5E79;	13'h1330: data <= 32'h5C66C441;	13'h1331: data <= 32'h5CA32A08;	13'h1332: data <= 32'h5CDF8FD0;	13'h1333: data <= 32'h5D1BF598;	13'h1334: data <= 32'h5D585B60;	13'h1335: data <= 32'h5D94C127;	13'h1336: data <= 32'h5DD126EF;	13'h1337: data <= 32'h5E0D8CB7;	13'h1338: data <= 32'h5E49F27E;	13'h1339: data <= 32'h5E865846;	13'h133A: data <= 32'h5EC2BE0E;	13'h133B: data <= 32'h5EFF23D5;	13'h133C: data <= 32'h5F3B899D;	13'h133D: data <= 32'h5F77EF65;	13'h133E: data <= 32'h5FB4552C;	13'h133F: data <= 32'h5FF0BAF4;	13'h1340: data <= 32'h602D20BC;	13'h1341: data <= 32'h60698684;	13'h1342: data <= 32'h60A5EC4B;	13'h1343: data <= 32'h60E25213;	13'h1344: data <= 32'h611EB7DB;	13'h1345: data <= 32'h615B1DA2;	13'h1346: data <= 32'h6197836A;	13'h1347: data <= 32'h61D3E932;	13'h1348: data <= 32'h62104EF9;	13'h1349: data <= 32'h624CB4C1;	13'h134A: data <= 32'h62891A89;	13'h134B: data <= 32'h62C58050;	13'h134C: data <= 32'h62FD02E2;	13'h134D: data <= 32'h6331582A;	13'h134E: data <= 32'h6365AD72;	13'h134F: data <= 32'h639A02BA;	13'h1350: data <= 32'h63CE5802;	13'h1351: data <= 32'h6402AD4A;	13'h1352: data <= 32'h64370292;	13'h1353: data <= 32'h646B57DA;	13'h1354: data <= 32'h649FAD22;	13'h1355: data <= 32'h64D4026A;	13'h1356: data <= 32'h650857B2;	13'h1357: data <= 32'h653CACFA;	13'h1358: data <= 32'h65710241;	13'h1359: data <= 32'h65A55789;	13'h135A: data <= 32'h65D9ACD1;	13'h135B: data <= 32'h660E0219;	13'h135C: data <= 32'h66425761;	13'h135D: data <= 32'h6676ACA9;	13'h135E: data <= 32'h66AB01F1;	13'h135F: data <= 32'h66DF5739;	13'h1360: data <= 32'h6713AC81;	13'h1361: data <= 32'h674801C9;	13'h1362: data <= 32'h677C5711;	13'h1363: data <= 32'h67B0AC59;	13'h1364: data <= 32'h67E501A1;	13'h1365: data <= 32'h681956E9;	13'h1366: data <= 32'h684DAC31;	13'h1367: data <= 32'h68820179;	13'h1368: data <= 32'h68B656C1;	13'h1369: data <= 32'h68EAAC09;	13'h136A: data <= 32'h691CD741;	13'h136B: data <= 32'h694A0823;	13'h136C: data <= 32'h69773905;	13'h136D: data <= 32'h69A469E6;	13'h136E: data <= 32'h69D19AC8;	13'h136F: data <= 32'h69FECBAA;	13'h1370: data <= 32'h6A2BFC8B;	13'h1371: data <= 32'h6A592D6D;	13'h1372: data <= 32'h6A865E4F;	13'h1373: data <= 32'h6AB38F30;	13'h1374: data <= 32'h6AE0C012;	13'h1375: data <= 32'h6B0DF0F4;	13'h1376: data <= 32'h6B3B21D5;	13'h1377: data <= 32'h6B6852B7;	13'h1378: data <= 32'h6B958399;	13'h1379: data <= 32'h6BC2B47A;	13'h137A: data <= 32'h6BEFE55C;	13'h137B: data <= 32'h6C1D163E;	13'h137C: data <= 32'h6C4A471F;	13'h137D: data <= 32'h6C777801;	13'h137E: data <= 32'h6CA4A8E3;	13'h137F: data <= 32'h6CD1D9C4;	13'h1380: data <= 32'h6CFF0AA6;	13'h1381: data <= 32'h6D2C3B88;	13'h1382: data <= 32'h6D596C69;	13'h1383: data <= 32'h6D869D4B;	13'h1384: data <= 32'h6DB3CE2D;	13'h1385: data <= 32'h6DE0FF0E;	13'h1386: data <= 32'h6E0E2FF0;	13'h1387: data <= 32'h6E3B60D2;	13'h1388: data <= 32'h6E6891B4;	13'h1389: data <= 32'h6E8FBBB3;	13'h138A: data <= 32'h6EB6E5B2;	13'h138B: data <= 32'h6EDE0FB2;	13'h138C: data <= 32'h6F0539B1;	13'h138D: data <= 32'h6F2C63B1;	13'h138E: data <= 32'h6F538DB0;	13'h138F: data <= 32'h6F7AB7B0;	13'h1390: data <= 32'h6FA1E1AF;	13'h1391: data <= 32'h6FC90BAF;	13'h1392: data <= 32'h6FF035AE;	13'h1393: data <= 32'h70175FAE;	13'h1394: data <= 32'h703E89AD;	13'h1395: data <= 32'h7065B3AD;	13'h1396: data <= 32'h708CDDAC;	13'h1397: data <= 32'h70B407AC;	13'h1398: data <= 32'h70DB31AB;	13'h1399: data <= 32'h71025BAB;	13'h139A: data <= 32'h712985AA;	13'h139B: data <= 32'h7150AFAA;	13'h139C: data <= 32'h7177D9A9;	13'h139D: data <= 32'h719F03A9;	13'h139E: data <= 32'h71C62DA8;	13'h139F: data <= 32'h71ED57A8;	13'h13A0: data <= 32'h721481A7;	13'h13A1: data <= 32'h723BABA7;	13'h13A2: data <= 32'h7262D5A6;	13'h13A3: data <= 32'h7289FFA6;	13'h13A4: data <= 32'h72B129A5;	13'h13A5: data <= 32'h72D853A5;	13'h13A6: data <= 32'h72FF7DA4;	13'h13A7: data <= 32'h7322CC50;	13'h13A8: data <= 32'h73446DB7;	13'h13A9: data <= 32'h73660F1D;	13'h13AA: data <= 32'h7387B084;	13'h13AB: data <= 32'h73A951EA;	13'h13AC: data <= 32'h73CAF351;	13'h13AD: data <= 32'h73EC94B7;	13'h13AE: data <= 32'h740E361E;	13'h13AF: data <= 32'h742FD784;	13'h13B0: data <= 32'h745178EA;	13'h13B1: data <= 32'h74731A51;	13'h13B2: data <= 32'h7494BBB7;	13'h13B3: data <= 32'h74B65D1E;	13'h13B4: data <= 32'h74D7FE84;	13'h13B5: data <= 32'h74F99FEB;	13'h13B6: data <= 32'h751B4151;	13'h13B7: data <= 32'h753CE2B8;	13'h13B8: data <= 32'h755E841E;	13'h13B9: data <= 32'h75802585;	13'h13BA: data <= 32'h75A1C6EB;	13'h13BB: data <= 32'h75C36852;	13'h13BC: data <= 32'h75E509B8;	13'h13BD: data <= 32'h7606AB1F;	13'h13BE: data <= 32'h76284C85;	13'h13BF: data <= 32'h7649EDEC;	13'h13C0: data <= 32'h766B8F52;	13'h13C1: data <= 32'h768D30B9;	13'h13C2: data <= 32'h76AED21F;	13'h13C3: data <= 32'h76D07386;	13'h13C4: data <= 32'h76F214EC;	13'h13C5: data <= 32'h771176F7;	13'h13C6: data <= 32'h772D63D7;	13'h13C7: data <= 32'h774950B8;	13'h13C8: data <= 32'h77653D98;	13'h13C9: data <= 32'h77812A79;	13'h13CA: data <= 32'h779D1759;	13'h13CB: data <= 32'h77B9043A;	13'h13CC: data <= 32'h77D4F11A;	13'h13CD: data <= 32'h77F0DDFB;	13'h13CE: data <= 32'h780CCADB;	13'h13CF: data <= 32'h7828B7BC;	13'h13D0: data <= 32'h7844A49C;	13'h13D1: data <= 32'h7860917D;	13'h13D2: data <= 32'h787C7E5D;	13'h13D3: data <= 32'h78986B3E;	13'h13D4: data <= 32'h78B4581E;	13'h13D5: data <= 32'h78D044FF;	13'h13D6: data <= 32'h78EC31DF;	13'h13D7: data <= 32'h79081EC0;	13'h13D8: data <= 32'h79240BA0;	13'h13D9: data <= 32'h793FF881;	13'h13DA: data <= 32'h795BE561;	13'h13DB: data <= 32'h7977D242;	13'h13DC: data <= 32'h7993BF22;	13'h13DD: data <= 32'h79AFAC02;	13'h13DE: data <= 32'h79CB98E3;	13'h13DF: data <= 32'h79E785C3;	13'h13E0: data <= 32'h7A0372A4;	13'h13E1: data <= 32'h7A1F5F84;	13'h13E2: data <= 32'h7A3B4C65;	13'h13E3: data <= 32'h7A56B280;	13'h13E4: data <= 32'h7A6CD4E4;	13'h13E5: data <= 32'h7A82F748;	13'h13E6: data <= 32'h7A9919AC;	13'h13E7: data <= 32'h7AAF3C10;	13'h13E8: data <= 32'h7AC55E74;	13'h13E9: data <= 32'h7ADB80D9;	13'h13EA: data <= 32'h7AF1A33D;	13'h13EB: data <= 32'h7B07C5A1;	13'h13EC: data <= 32'h7B1DE805;	13'h13ED: data <= 32'h7B340A69;	13'h13EE: data <= 32'h7B4A2CCD;	13'h13EF: data <= 32'h7B604F31;	13'h13F0: data <= 32'h7B767195;	13'h13F1: data <= 32'h7B8C93F9;	13'h13F2: data <= 32'h7BA2B65E;	13'h13F3: data <= 32'h7BB8D8C2;	13'h13F4: data <= 32'h7BCEFB26;	13'h13F5: data <= 32'h7BE51D8A;	13'h13F6: data <= 32'h7BFB3FEE;	13'h13F7: data <= 32'h7C116252;	13'h13F8: data <= 32'h7C2784B6;	13'h13F9: data <= 32'h7C3DA71A;	13'h13FA: data <= 32'h7C53C97E;	13'h13FB: data <= 32'h7C69EBE3;	13'h13FC: data <= 32'h7C800E47;	13'h13FD: data <= 32'h7C9630AB;	13'h13FE: data <= 32'h7CAC530F;	13'h13FF: data <= 32'h7CC27573;	13'h1400: data <= 32'h7CD897D7;	13'h1401: data <= 32'h7CEEBA3B;	13'h1402: data <= 32'h7D002158;	13'h1403: data <= 32'h7D104257;	13'h1404: data <= 32'h7D206357;	13'h1405: data <= 32'h7D308456;	13'h1406: data <= 32'h7D40A556;	13'h1407: data <= 32'h7D50C655;	13'h1408: data <= 32'h7D60E755;	13'h1409: data <= 32'h7D710854;	13'h140A: data <= 32'h7D812954;	13'h140B: data <= 32'h7D914A53;	13'h140C: data <= 32'h7DA16B53;	13'h140D: data <= 32'h7DB18C52;	13'h140E: data <= 32'h7DC1AD52;	13'h140F: data <= 32'h7DD1CE51;	13'h1410: data <= 32'h7DE1EF51;	13'h1411: data <= 32'h7DF21050;	13'h1412: data <= 32'h7E023150;	13'h1413: data <= 32'h7E12524F;	13'h1414: data <= 32'h7E22734F;	13'h1415: data <= 32'h7E32944E;	13'h1416: data <= 32'h7E42B54E;	13'h1417: data <= 32'h7E52D64D;	13'h1418: data <= 32'h7E62F74D;	13'h1419: data <= 32'h7E73184C;	13'h141A: data <= 32'h7E83394C;	13'h141B: data <= 32'h7E935A4B;	13'h141C: data <= 32'h7EA37B4B;	13'h141D: data <= 32'h7EB39C4A;	13'h141E: data <= 32'h7EC3BD4A;	13'h141F: data <= 32'h7ED3DE49;	13'h1420: data <= 32'h7EE09E16;	13'h1421: data <= 32'h7EE9C69C;	13'h1422: data <= 32'h7EF2EF22;	13'h1423: data <= 32'h7EFC17A8;	13'h1424: data <= 32'h7F05402E;	13'h1425: data <= 32'h7F0E68B5;	13'h1426: data <= 32'h7F17913B;	13'h1427: data <= 32'h7F20B9C1;	13'h1428: data <= 32'h7F29E247;	13'h1429: data <= 32'h7F330ACD;	13'h142A: data <= 32'h7F3C3354;	13'h142B: data <= 32'h7F455BDA;	13'h142C: data <= 32'h7F4E8460;	13'h142D: data <= 32'h7F57ACE6;	13'h142E: data <= 32'h7F60D56C;	13'h142F: data <= 32'h7F69FDF3;	13'h1430: data <= 32'h7F732679;	13'h1431: data <= 32'h7F7C4EFF;	13'h1432: data <= 32'h7F857785;	13'h1433: data <= 32'h7F8EA00B;	13'h1434: data <= 32'h7F97C892;	13'h1435: data <= 32'h7FA0F118;	13'h1436: data <= 32'h7FAA199E;	13'h1437: data <= 32'h7FB34224;	13'h1438: data <= 32'h7FBC6AAA;	13'h1439: data <= 32'h7FC59330;	13'h143A: data <= 32'h7FCEBBB7;	13'h143B: data <= 32'h7FD7E43D;	13'h143C: data <= 32'h7FE10CC3;	13'h143D: data <= 32'h7FEA3549;	13'h143E: data <= 32'h7FF1C97F;	13'h143F: data <= 32'h7FF2424B;	13'h1440: data <= 32'h7FF2BB16;	13'h1441: data <= 32'h7FF333E2;	13'h1442: data <= 32'h7FF3ACAD;	13'h1443: data <= 32'h7FF42579;	13'h1444: data <= 32'h7FF49E44;	13'h1445: data <= 32'h7FF51710;	13'h1446: data <= 32'h7FF58FDC;	13'h1447: data <= 32'h7FF608A7;	13'h1448: data <= 32'h7FF68173;	13'h1449: data <= 32'h7FF6FA3E;	13'h144A: data <= 32'h7FF7730A;	13'h144B: data <= 32'h7FF7EBD5;	13'h144C: data <= 32'h7FF864A1;	13'h144D: data <= 32'h7FF8DD6D;	13'h144E: data <= 32'h7FF95638;	13'h144F: data <= 32'h7FF9CF04;	13'h1450: data <= 32'h7FFA47CF;	13'h1451: data <= 32'h7FFAC09B;	13'h1452: data <= 32'h7FFB3966;	13'h1453: data <= 32'h7FFBB232;	13'h1454: data <= 32'h7FFC2AFE;	13'h1455: data <= 32'h7FFCA3C9;	13'h1456: data <= 32'h7FFD1C95;	13'h1457: data <= 32'h7FFD9560;	13'h1458: data <= 32'h7FFE0E2C;	13'h1459: data <= 32'h7FFE86F7;	13'h145A: data <= 32'h7FFEFFC3;	13'h145B: data <= 32'h7FFF788F;	13'h145C: data <= 32'h7FFFF15A;	13'h145D: data <= 32'h7FF72900;	13'h145E: data <= 32'h7FED19DD;	13'h145F: data <= 32'h7FE30ABB;	13'h1460: data <= 32'h7FD8FB99;	13'h1461: data <= 32'h7FCEEC77;	13'h1462: data <= 32'h7FC4DD55;	13'h1463: data <= 32'h7FBACE33;	13'h1464: data <= 32'h7FB0BF11;	13'h1465: data <= 32'h7FA6AFEF;	13'h1466: data <= 32'h7F9CA0CD;	13'h1467: data <= 32'h7F9291AB;	13'h1468: data <= 32'h7F888288;	13'h1469: data <= 32'h7F7E7366;	13'h146A: data <= 32'h7F746444;	13'h146B: data <= 32'h7F6A5522;	13'h146C: data <= 32'h7F604600;	13'h146D: data <= 32'h7F5636DE;	13'h146E: data <= 32'h7F4C27BC;	13'h146F: data <= 32'h7F42189A;	13'h1470: data <= 32'h7F380978;	13'h1471: data <= 32'h7F2DFA56;	13'h1472: data <= 32'h7F23EB33;	13'h1473: data <= 32'h7F19DC11;	13'h1474: data <= 32'h7F0FCCEF;	13'h1475: data <= 32'h7F05BDCD;	13'h1476: data <= 32'h7EFBAEAB;	13'h1477: data <= 32'h7EF19F89;	13'h1478: data <= 32'h7EE79067;	13'h1479: data <= 32'h7EDD8145;	13'h147A: data <= 32'h7ED37223;	13'h147B: data <= 32'h7EC25C38;	13'h147C: data <= 32'h7EAC18E2;	13'h147D: data <= 32'h7E95D58C;	13'h147E: data <= 32'h7E7F9237;	13'h147F: data <= 32'h7E694EE1;	13'h1480: data <= 32'h7E530B8B;	13'h1481: data <= 32'h7E3CC835;	13'h1482: data <= 32'h7E2684E0;	13'h1483: data <= 32'h7E10418A;	13'h1484: data <= 32'h7DF9FE34;	13'h1485: data <= 32'h7DE3BADE;	13'h1486: data <= 32'h7DCD7788;	13'h1487: data <= 32'h7DB73433;	13'h1488: data <= 32'h7DA0F0DD;	13'h1489: data <= 32'h7D8AAD87;	13'h148A: data <= 32'h7D746A31;	13'h148B: data <= 32'h7D5E26DB;	13'h148C: data <= 32'h7D47E386;	13'h148D: data <= 32'h7D31A030;	13'h148E: data <= 32'h7D1B5CDA;	13'h148F: data <= 32'h7D051984;	13'h1490: data <= 32'h7CEED62E;	13'h1491: data <= 32'h7CD892D9;	13'h1492: data <= 32'h7CC24F83;	13'h1493: data <= 32'h7CAC0C2D;	13'h1494: data <= 32'h7C95C8D7;	13'h1495: data <= 32'h7C7F8581;	13'h1496: data <= 32'h7C69422C;	13'h1497: data <= 32'h7C52FED6;	13'h1498: data <= 32'h7C3CBB80;	13'h1499: data <= 32'h7C22C2C6;	13'h149A: data <= 32'h7BFEE658;	13'h149B: data <= 32'h7BDB09E9;	13'h149C: data <= 32'h7BB72D7B;	13'h149D: data <= 32'h7B93510C;	13'h149E: data <= 32'h7B6F749E;	13'h149F: data <= 32'h7B4B982F;	13'h14A0: data <= 32'h7B27BBC1;	13'h14A1: data <= 32'h7B03DF52;	13'h14A2: data <= 32'h7AE002E4;	13'h14A3: data <= 32'h7ABC2675;	13'h14A4: data <= 32'h7A984A07;	13'h14A5: data <= 32'h7A746D98;	13'h14A6: data <= 32'h7A509129;	13'h14A7: data <= 32'h7A2CB4BB;	13'h14A8: data <= 32'h7A08D84C;	13'h14A9: data <= 32'h79E4FBDE;	13'h14AA: data <= 32'h79C11F6F;	13'h14AB: data <= 32'h799D4301;	13'h14AC: data <= 32'h79796692;	13'h14AD: data <= 32'h79558A24;	13'h14AE: data <= 32'h7931ADB5;	13'h14AF: data <= 32'h790DD147;	13'h14B0: data <= 32'h78E9F4D8;	13'h14B1: data <= 32'h78C6186A;	13'h14B2: data <= 32'h78A23BFB;	13'h14B3: data <= 32'h787E5F8D;	13'h14B4: data <= 32'h785A831E;	13'h14B5: data <= 32'h7836A6AF;	13'h14B6: data <= 32'h7812CA41;	13'h14B7: data <= 32'h77EEEDD2;	13'h14B8: data <= 32'h77BDAC8A;	13'h14B9: data <= 32'h778C001A;	13'h14BA: data <= 32'h775A53AB;	13'h14BB: data <= 32'h7728A73B;	13'h14BC: data <= 32'h76F6FACC;	13'h14BD: data <= 32'h76C54E5C;	13'h14BE: data <= 32'h7693A1ED;	13'h14BF: data <= 32'h7661F57D;	13'h14C0: data <= 32'h7630490D;	13'h14C1: data <= 32'h75FE9C9E;	13'h14C2: data <= 32'h75CCF02E;	13'h14C3: data <= 32'h759B43BF;	13'h14C4: data <= 32'h7569974F;	13'h14C5: data <= 32'h7537EAE0;	13'h14C6: data <= 32'h75063E70;	13'h14C7: data <= 32'h74D49201;	13'h14C8: data <= 32'h74A2E591;	13'h14C9: data <= 32'h74713922;	13'h14CA: data <= 32'h743F8CB2;	13'h14CB: data <= 32'h740DE043;	13'h14CC: data <= 32'h73DC33D3;	13'h14CD: data <= 32'h73AA8764;	13'h14CE: data <= 32'h7378DAF4;	13'h14CF: data <= 32'h73472E85;	13'h14D0: data <= 32'h73158215;	13'h14D1: data <= 32'h72E3D5A5;	13'h14D2: data <= 32'h72B22936;	13'h14D3: data <= 32'h72807CC6;	13'h14D4: data <= 32'h724ED057;	13'h14D5: data <= 32'h721D23E7;	13'h14D6: data <= 32'h71E2C992;	13'h14D7: data <= 32'h71A41849;	13'h14D8: data <= 32'h71656701;	13'h14D9: data <= 32'h7126B5B8;	13'h14DA: data <= 32'h70E8046F;	13'h14DB: data <= 32'h70A95327;	13'h14DC: data <= 32'h706AA1DE;	13'h14DD: data <= 32'h702BF095;	13'h14DE: data <= 32'h6FED3F4D;	13'h14DF: data <= 32'h6FAE8E04;	13'h14E0: data <= 32'h6F6FDCBC;	13'h14E1: data <= 32'h6F312B73;	13'h14E2: data <= 32'h6EF27A2A;	13'h14E3: data <= 32'h6EB3C8E2;	13'h14E4: data <= 32'h6E751799;	13'h14E5: data <= 32'h6E366650;	13'h14E6: data <= 32'h6DF7B508;	13'h14E7: data <= 32'h6DB903BF;	13'h14E8: data <= 32'h6D7A5277;	13'h14E9: data <= 32'h6D3BA12E;	13'h14EA: data <= 32'h6CFCEFE5;	13'h14EB: data <= 32'h6CBE3E9D;	13'h14EC: data <= 32'h6C7F8D54;	13'h14ED: data <= 32'h6C40DC0B;	13'h14EE: data <= 32'h6C022AC3;	13'h14EF: data <= 32'h6BC3797A;	13'h14F0: data <= 32'h6B84C832;	13'h14F1: data <= 32'h6B4616E9;	13'h14F2: data <= 32'h6B0765A0;	13'h14F3: data <= 32'h6AC8B458;	13'h14F4: data <= 32'h6A85DEDB;	13'h14F5: data <= 32'h6A3BCA04;	13'h14F6: data <= 32'h69F1B52D;	13'h14F7: data <= 32'h69A7A057;	13'h14F8: data <= 32'h695D8B80;	13'h14F9: data <= 32'h691376A9;	13'h14FA: data <= 32'h68C961D2;	13'h14FB: data <= 32'h687F4CFB;	13'h14FC: data <= 32'h68353824;	13'h14FD: data <= 32'h67EB234D;	13'h14FE: data <= 32'h67A10E76;	13'h14FF: data <= 32'h6756F99F;	13'h1500: data <= 32'h670CE4C8;	13'h1501: data <= 32'h66C2CFF1;	13'h1502: data <= 32'h6678BB1A;	13'h1503: data <= 32'h662EA643;	13'h1504: data <= 32'h65E4916C;	13'h1505: data <= 32'h659A7C95;	13'h1506: data <= 32'h655067BE;	13'h1507: data <= 32'h650652E7;	13'h1508: data <= 32'h64BC3E11;	13'h1509: data <= 32'h6472293A;	13'h150A: data <= 32'h64281463;	13'h150B: data <= 32'h63DDFF8C;	13'h150C: data <= 32'h6393EAB5;	13'h150D: data <= 32'h6349D5DE;	13'h150E: data <= 32'h62FFC107;	13'h150F: data <= 32'h62B5AC30;	13'h1510: data <= 32'h626B9759;	13'h1511: data <= 32'h62218282;	13'h1512: data <= 32'h61D6E8E5;	13'h1513: data <= 32'h61844545;	13'h1514: data <= 32'h6131A1A5;	13'h1515: data <= 32'h60DEFE05;	13'h1516: data <= 32'h608C5A65;	13'h1517: data <= 32'h6039B6C6;	13'h1518: data <= 32'h5FE71326;	13'h1519: data <= 32'h5F946F86;	13'h151A: data <= 32'h5F41CBE6;	13'h151B: data <= 32'h5EEF2846;	13'h151C: data <= 32'h5E9C84A6;	13'h151D: data <= 32'h5E49E106;	13'h151E: data <= 32'h5DF73D67;	13'h151F: data <= 32'h5DA499C7;	13'h1520: data <= 32'h5D51F627;	13'h1521: data <= 32'h5CFF5287;	13'h1522: data <= 32'h5CACAEE7;	13'h1523: data <= 32'h5C5A0B47;	13'h1524: data <= 32'h5C0767A8;	13'h1525: data <= 32'h5BB4C408;	13'h1526: data <= 32'h5B622068;	13'h1527: data <= 32'h5B0F7CC8;	13'h1528: data <= 32'h5ABCD928;	13'h1529: data <= 32'h5A6A3588;	13'h152A: data <= 32'h5A1791E8;	13'h152B: data <= 32'h59C4EE49;	13'h152C: data <= 32'h59724AA9;	13'h152D: data <= 32'h591FA709;	13'h152E: data <= 32'h58CD0369;	13'h152F: data <= 32'h587A5FC9;	13'h1530: data <= 32'h5827BC29;	13'h1531: data <= 32'h57D1D04C;	13'h1532: data <= 32'h577AD78D;	13'h1533: data <= 32'h5723DECF;	13'h1534: data <= 32'h56CCE610;	13'h1535: data <= 32'h5675ED52;	13'h1536: data <= 32'h561EF494;	13'h1537: data <= 32'h55C7FBD5;	13'h1538: data <= 32'h55710317;	13'h1539: data <= 32'h551A0A58;	13'h153A: data <= 32'h54C3119A;	13'h153B: data <= 32'h546C18DC;	13'h153C: data <= 32'h5415201D;	13'h153D: data <= 32'h53BE275F;	13'h153E: data <= 32'h53672EA1;	13'h153F: data <= 32'h531035E2;	13'h1540: data <= 32'h52B93D24;	13'h1541: data <= 32'h52624465;	13'h1542: data <= 32'h520B4BA7;	13'h1543: data <= 32'h51B452E9;	13'h1544: data <= 32'h515D5A2A;	13'h1545: data <= 32'h5106616C;	13'h1546: data <= 32'h50AF68AD;	13'h1547: data <= 32'h50586FEF;	13'h1548: data <= 32'h50017731;	13'h1549: data <= 32'h4FAA7E72;	13'h154A: data <= 32'h4F5385B4;	13'h154B: data <= 32'h4EFC8CF6;	13'h154C: data <= 32'h4EA59437;	13'h154D: data <= 32'h4E4E9B79;	13'h154E: data <= 32'h4DF7A2BA;	13'h154F: data <= 32'h4DA0A9FC;	13'h1550: data <= 32'h4D49B13E;	13'h1551: data <= 32'h4CF2B87F;	13'h1552: data <= 32'h4C9BBFC1;	13'h1553: data <= 32'h4C44C703;	13'h1554: data <= 32'h4BEDCE44;	13'h1555: data <= 32'h4B96D586;	13'h1556: data <= 32'h4B3FDCC7;	13'h1557: data <= 32'h4AE8E409;	13'h1558: data <= 32'h4A91EB4B;	13'h1559: data <= 32'h4A3AF28C;	13'h155A: data <= 32'h49E3F9CE;	13'h155B: data <= 32'h498D0110;	13'h155C: data <= 32'h49360851;	13'h155D: data <= 32'h48DF0F93;	13'h155E: data <= 32'h488816D5;	13'h155F: data <= 32'h48311E16;	13'h1560: data <= 32'h47DA2558;	13'h1561: data <= 32'h47832C9A;	13'h1562: data <= 32'h472C33DB;	13'h1563: data <= 32'h46D53B1D;	13'h1564: data <= 32'h467E425F;	13'h1565: data <= 32'h462749A0;	13'h1566: data <= 32'h45D050E2;	13'h1567: data <= 32'h45795823;	13'h1568: data <= 32'h45225F65;	13'h1569: data <= 32'h44CB66A7;	13'h156A: data <= 32'h44746DE8;	13'h156B: data <= 32'h441D752A;	13'h156C: data <= 32'h43C67C6C;	13'h156D: data <= 32'h43702293;	13'h156E: data <= 32'h431D428D;	13'h156F: data <= 32'h42CA6288;	13'h1570: data <= 32'h42778282;	13'h1571: data <= 32'h4224A27C;	13'h1572: data <= 32'h41D1C277;	13'h1573: data <= 32'h417EE271;	13'h1574: data <= 32'h412C026C;	13'h1575: data <= 32'h40D92266;	13'h1576: data <= 32'h40864260;	13'h1577: data <= 32'h4033625B;	13'h1578: data <= 32'h3FE08255;	13'h1579: data <= 32'h3F8DA24F;	13'h157A: data <= 32'h3F3AC24A;	13'h157B: data <= 32'h3EE7E244;	13'h157C: data <= 32'h3E95023F;	13'h157D: data <= 32'h3E422239;	13'h157E: data <= 32'h3DEF4233;	13'h157F: data <= 32'h3D9C622E;	13'h1580: data <= 32'h3D498228;	13'h1581: data <= 32'h3CF6A222;	13'h1582: data <= 32'h3CA3C21D;	13'h1583: data <= 32'h3C50E217;	13'h1584: data <= 32'h3BFE0211;	13'h1585: data <= 32'h3BAB220C;	13'h1586: data <= 32'h3B584206;	13'h1587: data <= 32'h3B056201;	13'h1588: data <= 32'h3AB281FB;	13'h1589: data <= 32'h3A5FA1F5;	13'h158A: data <= 32'h3A0CC1F0;	13'h158B: data <= 32'h39B9E1EA;	13'h158C: data <= 32'h396DE2E8;	13'h158D: data <= 32'h39231E5D;	13'h158E: data <= 32'h38D859D3;	13'h158F: data <= 32'h388D9548;	13'h1590: data <= 32'h3842D0BD;	13'h1591: data <= 32'h37F80C33;	13'h1592: data <= 32'h37AD47A8;	13'h1593: data <= 32'h3762831D;	13'h1594: data <= 32'h3717BE93;	13'h1595: data <= 32'h36CCFA08;	13'h1596: data <= 32'h3682357D;	13'h1597: data <= 32'h363770F3;	13'h1598: data <= 32'h35ECAC68;	13'h1599: data <= 32'h35A1E7DD;	13'h159A: data <= 32'h35572353;	13'h159B: data <= 32'h350C5EC8;	13'h159C: data <= 32'h34C19A3D;	13'h159D: data <= 32'h3476D5B3;	13'h159E: data <= 32'h342C1128;	13'h159F: data <= 32'h33E14C9D;	13'h15A0: data <= 32'h33968813;	13'h15A1: data <= 32'h334BC388;	13'h15A2: data <= 32'h3300FEFD;	13'h15A3: data <= 32'h32B63A73;	13'h15A4: data <= 32'h326B75E8;	13'h15A5: data <= 32'h3220B15D;	13'h15A6: data <= 32'h31D5ECD3;	13'h15A7: data <= 32'h318B2848;	13'h15A8: data <= 32'h314063BD;	13'h15A9: data <= 32'h30F59F33;	13'h15AA: data <= 32'h30B116F3;	13'h15AB: data <= 32'h3071C0F2;	13'h15AC: data <= 32'h30326AF1;	13'h15AD: data <= 32'h2FF314F0;	13'h15AE: data <= 32'h2FB3BEEE;	13'h15AF: data <= 32'h2F7468ED;	13'h15B0: data <= 32'h2F3512EC;	13'h15B1: data <= 32'h2EF5BCEB;	13'h15B2: data <= 32'h2EB666EA;	13'h15B3: data <= 32'h2E7710E9;	13'h15B4: data <= 32'h2E37BAE8;	13'h15B5: data <= 32'h2DF864E7;	13'h15B6: data <= 32'h2DB90EE6;	13'h15B7: data <= 32'h2D79B8E4;	13'h15B8: data <= 32'h2D3A62E3;	13'h15B9: data <= 32'h2CFB0CE2;	13'h15BA: data <= 32'h2CBBB6E1;	13'h15BB: data <= 32'h2C7C60E0;	13'h15BC: data <= 32'h2C3D0ADF;	13'h15BD: data <= 32'h2BFDB4DE;	13'h15BE: data <= 32'h2BBE5EDD;	13'h15BF: data <= 32'h2B7F08DC;	13'h15C0: data <= 32'h2B3FB2DA;	13'h15C1: data <= 32'h2B005CD9;	13'h15C2: data <= 32'h2AC106D8;	13'h15C3: data <= 32'h2A81B0D7;	13'h15C4: data <= 32'h2A425AD6;	13'h15C5: data <= 32'h2A0304D5;	13'h15C6: data <= 32'h29C3AED4;	13'h15C7: data <= 32'h298458D3;	13'h15C8: data <= 32'h2948500D;	13'h15C9: data <= 32'h291698A3;	13'h15CA: data <= 32'h28E4E138;	13'h15CB: data <= 32'h28B329CD;	13'h15CC: data <= 32'h28817262;	13'h15CD: data <= 32'h284FBAF7;	13'h15CE: data <= 32'h281E038D;	13'h15CF: data <= 32'h27EC4C22;	13'h15D0: data <= 32'h27BA94B7;	13'h15D1: data <= 32'h2788DD4C;	13'h15D2: data <= 32'h275725E2;	13'h15D3: data <= 32'h27256E77;	13'h15D4: data <= 32'h26F3B70C;	13'h15D5: data <= 32'h26C1FFA1;	13'h15D6: data <= 32'h26904837;	13'h15D7: data <= 32'h265E90CC;	13'h15D8: data <= 32'h262CD961;	13'h15D9: data <= 32'h25FB21F6;	13'h15DA: data <= 32'h25C96A8B;	13'h15DB: data <= 32'h2597B321;	13'h15DC: data <= 32'h2565FBB6;	13'h15DD: data <= 32'h2534444B;	13'h15DE: data <= 32'h25028CE0;	13'h15DF: data <= 32'h24D0D576;	13'h15E0: data <= 32'h249F1E0B;	13'h15E1: data <= 32'h246D66A0;	13'h15E2: data <= 32'h243BAF35;	13'h15E3: data <= 32'h2409F7CB;	13'h15E4: data <= 32'h23D84060;	13'h15E5: data <= 32'h23A688F5;	13'h15E6: data <= 32'h2374D18A;	13'h15E7: data <= 32'h23512F82;	13'h15E8: data <= 32'h232E7616;	13'h15E9: data <= 32'h230BBCA9;	13'h15EA: data <= 32'h22E9033C;	13'h15EB: data <= 32'h22C649CF;	13'h15EC: data <= 32'h22A39062;	13'h15ED: data <= 32'h2280D6F5;	13'h15EE: data <= 32'h225E1D88;	13'h15EF: data <= 32'h223B641B;	13'h15F0: data <= 32'h2218AAAF;	13'h15F1: data <= 32'h21F5F142;	13'h15F2: data <= 32'h21D337D5;	13'h15F3: data <= 32'h21B07E68;	13'h15F4: data <= 32'h218DC4FB;	13'h15F5: data <= 32'h216B0B8E;	13'h15F6: data <= 32'h21485221;	13'h15F7: data <= 32'h212598B4;	13'h15F8: data <= 32'h2102DF48;	13'h15F9: data <= 32'h20E025DB;	13'h15FA: data <= 32'h20BD6C6E;	13'h15FB: data <= 32'h209AB301;	13'h15FC: data <= 32'h2077F994;	13'h15FD: data <= 32'h20554027;	13'h15FE: data <= 32'h203286BA;	13'h15FF: data <= 32'h200FCD4E;	13'h1600: data <= 32'h1FED13E1;	13'h1601: data <= 32'h1FCA5A74;	13'h1602: data <= 32'h1FA7A107;	13'h1603: data <= 32'h1F84E79A;	13'h1604: data <= 32'h1F622E2D;	13'h1605: data <= 32'h1F48E6A7;	13'h1606: data <= 32'h1F3504C8;	13'h1607: data <= 32'h1F2122EA;	13'h1608: data <= 32'h1F0D410B;	13'h1609: data <= 32'h1EF95F2D;	13'h160A: data <= 32'h1EE57D4F;	13'h160B: data <= 32'h1ED19B70;	13'h160C: data <= 32'h1EBDB992;	13'h160D: data <= 32'h1EA9D7B4;	13'h160E: data <= 32'h1E95F5D5;	13'h160F: data <= 32'h1E8213F7;	13'h1610: data <= 32'h1E6E3218;	13'h1611: data <= 32'h1E5A503A;	13'h1612: data <= 32'h1E466E5C;	13'h1613: data <= 32'h1E328C7D;	13'h1614: data <= 32'h1E1EAA9F;	13'h1615: data <= 32'h1E0AC8C0;	13'h1616: data <= 32'h1DF6E6E2;	13'h1617: data <= 32'h1DE30504;	13'h1618: data <= 32'h1DCF2325;	13'h1619: data <= 32'h1DBB4147;	13'h161A: data <= 32'h1DA75F69;	13'h161B: data <= 32'h1D937D8A;	13'h161C: data <= 32'h1D7F9BAC;	13'h161D: data <= 32'h1D6BB9CD;	13'h161E: data <= 32'h1D57D7EF;	13'h161F: data <= 32'h1D43F611;	13'h1620: data <= 32'h1D301432;	13'h1621: data <= 32'h1D1C3254;	13'h1622: data <= 32'h1D085075;	13'h1623: data <= 32'h1CF88EA2;	13'h1624: data <= 32'h1CF10CE4;	13'h1625: data <= 32'h1CE98B26;	13'h1626: data <= 32'h1CE20969;	13'h1627: data <= 32'h1CDA87AB;	13'h1628: data <= 32'h1CD305ED;	13'h1629: data <= 32'h1CCB8430;	13'h162A: data <= 32'h1CC40272;	13'h162B: data <= 32'h1CBC80B4;	13'h162C: data <= 32'h1CB4FEF6;	13'h162D: data <= 32'h1CAD7D39;	13'h162E: data <= 32'h1CA5FB7B;	13'h162F: data <= 32'h1C9E79BD;	13'h1630: data <= 32'h1C96F800;	13'h1631: data <= 32'h1C8F7642;	13'h1632: data <= 32'h1C87F484;	13'h1633: data <= 32'h1C8072C6;	13'h1634: data <= 32'h1C78F109;	13'h1635: data <= 32'h1C716F4B;	13'h1636: data <= 32'h1C69ED8D;	13'h1637: data <= 32'h1C626BD0;	13'h1638: data <= 32'h1C5AEA12;	13'h1639: data <= 32'h1C536854;	13'h163A: data <= 32'h1C4BE696;	13'h163B: data <= 32'h1C4464D9;	13'h163C: data <= 32'h1C3CE31B;	13'h163D: data <= 32'h1C35615D;	13'h163E: data <= 32'h1C2DDFA0;	13'h163F: data <= 32'h1C265DE2;	13'h1640: data <= 32'h1C1EDC24;	13'h1641: data <= 32'h1C1799A0;	13'h1642: data <= 32'h1C183E59;	13'h1643: data <= 32'h1C18E311;	13'h1644: data <= 32'h1C1987CA;	13'h1645: data <= 32'h1C1A2C82;	13'h1646: data <= 32'h1C1AD13B;	13'h1647: data <= 32'h1C1B75F3;	13'h1648: data <= 32'h1C1C1AAC;	13'h1649: data <= 32'h1C1CBF64;	13'h164A: data <= 32'h1C1D641D;	13'h164B: data <= 32'h1C1E08D5;	13'h164C: data <= 32'h1C1EAD8E;	13'h164D: data <= 32'h1C1F5246;	13'h164E: data <= 32'h1C1FF6FF;	13'h164F: data <= 32'h1C209BB7;	13'h1650: data <= 32'h1C214070;	13'h1651: data <= 32'h1C21E528;	13'h1652: data <= 32'h1C2289E1;	13'h1653: data <= 32'h1C232E99;	13'h1654: data <= 32'h1C23D352;	13'h1655: data <= 32'h1C24780A;	13'h1656: data <= 32'h1C251CC3;	13'h1657: data <= 32'h1C25C17B;	13'h1658: data <= 32'h1C266634;	13'h1659: data <= 32'h1C270AEC;	13'h165A: data <= 32'h1C27AFA5;	13'h165B: data <= 32'h1C28545D;	13'h165C: data <= 32'h1C28F916;	13'h165D: data <= 32'h1C299DCE;	13'h165E: data <= 32'h1C2A4287;	13'h165F: data <= 32'h1C2AE73F;	13'h1660: data <= 32'h1C2E2ED3;	13'h1661: data <= 32'h1C327378;	13'h1662: data <= 32'h1C36B81E;	13'h1663: data <= 32'h1C3AFCC3;	13'h1664: data <= 32'h1C3F4169;	13'h1665: data <= 32'h1C43860F;	13'h1666: data <= 32'h1C47CAB4;	13'h1667: data <= 32'h1C4C0F5A;	13'h1668: data <= 32'h1C505400;	13'h1669: data <= 32'h1C5498A5;	13'h166A: data <= 32'h1C58DD4B;	13'h166B: data <= 32'h1C5D21F1;	13'h166C: data <= 32'h1C616696;	13'h166D: data <= 32'h1C65AB3C;	13'h166E: data <= 32'h1C69EFE1;	13'h166F: data <= 32'h1C6E3487;	13'h1670: data <= 32'h1C72792D;	13'h1671: data <= 32'h1C76BDD2;	13'h1672: data <= 32'h1C7B0278;	13'h1673: data <= 32'h1C7F471E;	13'h1674: data <= 32'h1C838BC3;	13'h1675: data <= 32'h1C87D069;	13'h1676: data <= 32'h1C8C150F;	13'h1677: data <= 32'h1C9059B4;	13'h1678: data <= 32'h1C949E5A;	13'h1679: data <= 32'h1C98E2FF;	13'h167A: data <= 32'h1C9D27A5;	13'h167B: data <= 32'h1CA16C4B;	13'h167C: data <= 32'h1CA5B0F0;	13'h167D: data <= 32'h1CA9F596;	13'h167E: data <= 32'h1CADBA1E;	13'h167F: data <= 32'h1CB0D0C7;	13'h1680: data <= 32'h1CB3E76F;	13'h1681: data <= 32'h1CB6FE18;	13'h1682: data <= 32'h1CBA14C1;	13'h1683: data <= 32'h1CBD2B6A;	13'h1684: data <= 32'h1CC04212;	13'h1685: data <= 32'h1CC358BB;	13'h1686: data <= 32'h1CC66F64;	13'h1687: data <= 32'h1CC9860D;	13'h1688: data <= 32'h1CCC9CB6;	13'h1689: data <= 32'h1CCFB35E;	13'h168A: data <= 32'h1CD2CA07;	13'h168B: data <= 32'h1CD5E0B0;	13'h168C: data <= 32'h1CD8F759;	13'h168D: data <= 32'h1CDC0E01;	13'h168E: data <= 32'h1CDF24AA;	13'h168F: data <= 32'h1CE23B53;	13'h1690: data <= 32'h1CE551FC;	13'h1691: data <= 32'h1CE868A4;	13'h1692: data <= 32'h1CEB7F4D;	13'h1693: data <= 32'h1CEE95F6;	13'h1694: data <= 32'h1CF1AC9F;	13'h1695: data <= 32'h1CF4C348;	13'h1696: data <= 32'h1CF7D9F0;	13'h1697: data <= 32'h1CFAF099;	13'h1698: data <= 32'h1CFE0742;	13'h1699: data <= 32'h1D011DEB;	13'h169A: data <= 32'h1D043493;	13'h169B: data <= 32'h1D074B3C;	13'h169C: data <= 32'h1D09A437;	13'h169D: data <= 32'h1D069E07;	13'h169E: data <= 32'h1D0397D7;	13'h169F: data <= 32'h1D0091A8;	13'h16A0: data <= 32'h1CFD8B78;	13'h16A1: data <= 32'h1CFA8548;	13'h16A2: data <= 32'h1CF77F18;	13'h16A3: data <= 32'h1CF478E8;	13'h16A4: data <= 32'h1CF172B8;	13'h16A5: data <= 32'h1CEE6C88;	13'h16A6: data <= 32'h1CEB6658;	13'h16A7: data <= 32'h1CE86028;	13'h16A8: data <= 32'h1CE559F9;	13'h16A9: data <= 32'h1CE253C9;	13'h16AA: data <= 32'h1CDF4D99;	13'h16AB: data <= 32'h1CDC4769;	13'h16AC: data <= 32'h1CD94139;	13'h16AD: data <= 32'h1CD63B09;	13'h16AE: data <= 32'h1CD334D9;	13'h16AF: data <= 32'h1CD02EA9;	13'h16B0: data <= 32'h1CCD2879;	13'h16B1: data <= 32'h1CCA2249;	13'h16B2: data <= 32'h1CC71C1A;	13'h16B3: data <= 32'h1CC415EA;	13'h16B4: data <= 32'h1CC10FBA;	13'h16B5: data <= 32'h1CBE098A;	13'h16B6: data <= 32'h1CBB035A;	13'h16B7: data <= 32'h1CB7FD2A;	13'h16B8: data <= 32'h1CB4F6FA;	13'h16B9: data <= 32'h1CB1F0CA;	13'h16BA: data <= 32'h1CAEEA9A;	13'h16BB: data <= 32'h1CA407D4;	13'h16BC: data <= 32'h1C9765D0;	13'h16BD: data <= 32'h1C8AC3CC;	13'h16BE: data <= 32'h1C7E21C8;	13'h16BF: data <= 32'h1C717FC4;	13'h16C0: data <= 32'h1C64DDC0;	13'h16C1: data <= 32'h1C583BBC;	13'h16C2: data <= 32'h1C4B99B8;	13'h16C3: data <= 32'h1C3EF7B4;	13'h16C4: data <= 32'h1C3255B0;	13'h16C5: data <= 32'h1C25B3AC;	13'h16C6: data <= 32'h1C1911A8;	13'h16C7: data <= 32'h1C0C6FA3;	13'h16C8: data <= 32'h1BFFCD9F;	13'h16C9: data <= 32'h1BF32B9B;	13'h16CA: data <= 32'h1BE68997;	13'h16CB: data <= 32'h1BD9E793;	13'h16CC: data <= 32'h1BCD458F;	13'h16CD: data <= 32'h1BC0A38B;	13'h16CE: data <= 32'h1BB40187;	13'h16CF: data <= 32'h1BA75F83;	13'h16D0: data <= 32'h1B9ABD7F;	13'h16D1: data <= 32'h1B8E1B7B;	13'h16D2: data <= 32'h1B817977;	13'h16D3: data <= 32'h1B74D773;	13'h16D4: data <= 32'h1B68356F;	13'h16D5: data <= 32'h1B5B936B;	13'h16D6: data <= 32'h1B4EF167;	13'h16D7: data <= 32'h1B424F63;	13'h16D8: data <= 32'h1B35AD5E;	13'h16D9: data <= 32'h1B235500;	13'h16DA: data <= 32'h1B0B9C4C;	13'h16DB: data <= 32'h1AF3E399;	13'h16DC: data <= 32'h1ADC2AE5;	13'h16DD: data <= 32'h1AC47231;	13'h16DE: data <= 32'h1AACB97E;	13'h16DF: data <= 32'h1A9500CA;	13'h16E0: data <= 32'h1A7D4816;	13'h16E1: data <= 32'h1A658F62;	13'h16E2: data <= 32'h1A4DD6AF;	13'h16E3: data <= 32'h1A361DFB;	13'h16E4: data <= 32'h1A1E6547;	13'h16E5: data <= 32'h1A06AC94;	13'h16E6: data <= 32'h19EEF3E0;	13'h16E7: data <= 32'h19D73B2C;	13'h16E8: data <= 32'h19BF8279;	13'h16E9: data <= 32'h19A7C9C5;	13'h16EA: data <= 32'h19901111;	13'h16EB: data <= 32'h1978585E;	13'h16EC: data <= 32'h19609FAA;	13'h16ED: data <= 32'h1948E6F6;	13'h16EE: data <= 32'h19312E43;	13'h16EF: data <= 32'h1919758F;	13'h16F0: data <= 32'h1901BCDB;	13'h16F1: data <= 32'h18EA0427;	13'h16F2: data <= 32'h18D24B74;	13'h16F3: data <= 32'h18BA92C0;	13'h16F4: data <= 32'h18A2DA0C;	13'h16F5: data <= 32'h188B2159;	13'h16F6: data <= 32'h187368A5;	13'h16F7: data <= 32'h1859432A;	13'h16F8: data <= 32'h18361BEC;	13'h16F9: data <= 32'h1812F4AF;	13'h16FA: data <= 32'h17EFCD72;	13'h16FB: data <= 32'h17CCA635;	13'h16FC: data <= 32'h17A97EF7;	13'h16FD: data <= 32'h178657BA;	13'h16FE: data <= 32'h1763307D;	13'h16FF: data <= 32'h17400940;	13'h1700: data <= 32'h171CE202;	13'h1701: data <= 32'h16F9BAC5;	13'h1702: data <= 32'h16D69388;	13'h1703: data <= 32'h16B36C4B;	13'h1704: data <= 32'h1690450D;	13'h1705: data <= 32'h166D1DD0;	13'h1706: data <= 32'h1649F693;	13'h1707: data <= 32'h1626CF56;	13'h1708: data <= 32'h1603A818;	13'h1709: data <= 32'h15E080DB;	13'h170A: data <= 32'h15BD599E;	13'h170B: data <= 32'h159A3261;	13'h170C: data <= 32'h15770B23;	13'h170D: data <= 32'h1553E3E6;	13'h170E: data <= 32'h1530BCA9;	13'h170F: data <= 32'h150D956C;	13'h1710: data <= 32'h14EA6E2F;	13'h1711: data <= 32'h14C746F1;	13'h1712: data <= 32'h14A41FB4;	13'h1713: data <= 32'h1480F877;	13'h1714: data <= 32'h145DD13A;	13'h1715: data <= 32'h143AA9FC;	13'h1716: data <= 32'h140DEAE9;	13'h1717: data <= 32'h13E03641;	13'h1718: data <= 32'h13B28198;	13'h1719: data <= 32'h1384CCF0;	13'h171A: data <= 32'h13571847;	13'h171B: data <= 32'h1329639F;	13'h171C: data <= 32'h12FBAEF6;	13'h171D: data <= 32'h12CDFA4E;	13'h171E: data <= 32'h12A045A5;	13'h171F: data <= 32'h127290FD;	13'h1720: data <= 32'h1244DC54;	13'h1721: data <= 32'h121727AC;	13'h1722: data <= 32'h11E97303;	13'h1723: data <= 32'h11BBBE5B;	13'h1724: data <= 32'h118E09B2;	13'h1725: data <= 32'h1160550A;	13'h1726: data <= 32'h1132A061;	13'h1727: data <= 32'h1104EBB9;	13'h1728: data <= 32'h10D73710;	13'h1729: data <= 32'h10A98268;	13'h172A: data <= 32'h107BCDC0;	13'h172B: data <= 32'h104E1917;	13'h172C: data <= 32'h1020646F;	13'h172D: data <= 32'h0FF2AFC6;	13'h172E: data <= 32'h0FC4FB1E;	13'h172F: data <= 32'h0F974675;	13'h1730: data <= 32'h0F6991CD;	13'h1731: data <= 32'h0F3BDD24;	13'h1732: data <= 32'h0F0E287C;	13'h1733: data <= 32'h0EE073D3;	13'h1734: data <= 32'h0EAE0A8B;	13'h1735: data <= 32'h0E789241;	13'h1736: data <= 32'h0E4319F8;	13'h1737: data <= 32'h0E0DA1AE;	13'h1738: data <= 32'h0DD82965;	13'h1739: data <= 32'h0DA2B11B;	13'h173A: data <= 32'h0D6D38D1;	13'h173B: data <= 32'h0D37C088;	13'h173C: data <= 32'h0D02483E;	13'h173D: data <= 32'h0CCCCFF5;	13'h173E: data <= 32'h0C9757AB;	13'h173F: data <= 32'h0C61DF61;	13'h1740: data <= 32'h0C2C6718;	13'h1741: data <= 32'h0BF6EECE;	13'h1742: data <= 32'h0BC17685;	13'h1743: data <= 32'h0B8BFE3B;	13'h1744: data <= 32'h0B5685F2;	13'h1745: data <= 32'h0B210DA8;	13'h1746: data <= 32'h0AEB955E;	13'h1747: data <= 32'h0AB61D15;	13'h1748: data <= 32'h0A80A4CB;	13'h1749: data <= 32'h0A4B2C82;	13'h174A: data <= 32'h0A15B438;	13'h174B: data <= 32'h09E03BEE;	13'h174C: data <= 32'h09AAC3A5;	13'h174D: data <= 32'h09754B5B;	13'h174E: data <= 32'h093FD312;	13'h174F: data <= 32'h090A5AC8;	13'h1750: data <= 32'h08D4E27E;	13'h1751: data <= 32'h089F6A35;	13'h1752: data <= 32'h0865CFB7;	13'h1753: data <= 32'h0822B359;	13'h1754: data <= 32'h07DF96FB;	13'h1755: data <= 32'h079C7A9E;	13'h1756: data <= 32'h07595E40;	13'h1757: data <= 32'h071641E3;	13'h1758: data <= 32'h06D32585;	13'h1759: data <= 32'h06900927;	13'h175A: data <= 32'h064CECCA;	13'h175B: data <= 32'h0609D06C;	13'h175C: data <= 32'h05C6B40F;	13'h175D: data <= 32'h058397B1;	13'h175E: data <= 32'h05407B53;	13'h175F: data <= 32'h04FD5EF6;	13'h1760: data <= 32'h04BA4298;	13'h1761: data <= 32'h0477263B;	13'h1762: data <= 32'h043409DD;	13'h1763: data <= 32'h03F0ED7F;	13'h1764: data <= 32'h03ADD122;	13'h1765: data <= 32'h036AB4C4;	13'h1766: data <= 32'h03279867;	13'h1767: data <= 32'h02E47C09;	13'h1768: data <= 32'h02A15FAB;	13'h1769: data <= 32'h025E434E;	13'h176A: data <= 32'h021B26F0;	13'h176B: data <= 32'h01D80A93;	13'h176C: data <= 32'h0194EE35;	13'h176D: data <= 32'h0151D1D7;	13'h176E: data <= 32'h010EB57A;	13'h176F: data <= 32'h00CB991C;endcase
    end
    endmodule