`timescale 1ns / 1ps
    module wave_rom (
    input clk,
    input en,
    input [13:0] addr,
    output reg [31:0] data
    );

    always @(posedge clk) begin
    if (en)
        case(addr)
			14'h0000: data <= 32'h00000000;	14'h0001: data <= 32'h0044A10B;	14'h0002: data <= 32'h00894204;	14'h0003: data <= 32'h00CDE2D4;	14'h0004: data <= 32'h0112836A;	14'h0005: data <= 32'h015723B1;	14'h0006: data <= 32'h019BC395;	14'h0007: data <= 32'h01E06302;	14'h0008: data <= 32'h022501E6;	14'h0009: data <= 32'h0269A02C;	14'h000A: data <= 32'h02AE3DC0;	14'h000B: data <= 32'h02F2DA8F;	14'h000C: data <= 32'h03377685;	14'h000D: data <= 32'h037C118E;	14'h000E: data <= 32'h03C0AB96;	14'h000F: data <= 32'h0405448B;	14'h0010: data <= 32'h0449DC58;	14'h0011: data <= 32'h048E72E9;	14'h0012: data <= 32'h04D3082A;	14'h0013: data <= 32'h05179C09;	14'h0014: data <= 32'h055C2E71;	14'h0015: data <= 32'h05A0BF4F;	14'h0016: data <= 32'h05E54E8E;	14'h0017: data <= 32'h0629DC1B;	14'h0018: data <= 32'h066E67E3;	14'h0019: data <= 32'h06B2F1D2;	14'h001A: data <= 32'h06F779D3;	14'h001B: data <= 32'h073BFFD4;	14'h001C: data <= 32'h078083C0;	14'h001D: data <= 32'h07C50585;	14'h001E: data <= 32'h0809850D;	14'h001F: data <= 32'h084E0246;	14'h0020: data <= 32'h08927D1C;	14'h0021: data <= 32'h08D6F57B;	14'h0022: data <= 32'h091B6B50;	14'h0023: data <= 32'h095FDE86;	14'h0024: data <= 32'h09A44F0B;	14'h0025: data <= 32'h09E8BCC9;	14'h0026: data <= 32'h0A2D27AF;	14'h0027: data <= 32'h0A718FA8;	14'h0028: data <= 32'h0AB5F4A0;	14'h0029: data <= 32'h0AFA5684;	14'h002A: data <= 32'h0B3EB53F;	14'h002B: data <= 32'h0B8310C0;	14'h002C: data <= 32'h0BC768F1;	14'h002D: data <= 32'h0C0BBDBF;	14'h002E: data <= 32'h0C500F17;	14'h002F: data <= 32'h0C945CE5;	14'h0030: data <= 32'h0CD8A715;	14'h0031: data <= 32'h0D1CED93;	14'h0032: data <= 32'h0D61304D;	14'h0033: data <= 32'h0DA56F2E;	14'h0034: data <= 32'h0DE9AA23;	14'h0035: data <= 32'h0E2DE117;	14'h0036: data <= 32'h0E7213F8;	14'h0037: data <= 32'h0EB642B3;	14'h0038: data <= 32'h0EFA6D32;	14'h0039: data <= 32'h0F3E9363;	14'h003A: data <= 32'h0F82B532;	14'h003B: data <= 32'h0FC6D28C;	14'h003C: data <= 32'h100AEB5D;	14'h003D: data <= 32'h104EFF91;	14'h003E: data <= 32'h10930F15;	14'h003F: data <= 32'h10D719D5;	14'h0040: data <= 32'h111B1FBE;	14'h0041: data <= 32'h115F20BC;	14'h0042: data <= 32'h11A31CBB;	14'h0043: data <= 32'h11E713A9;	14'h0044: data <= 32'h122B0571;	14'h0045: data <= 32'h126EF200;	14'h0046: data <= 32'h12B2D942;	14'h0047: data <= 32'h12F6BB25;	14'h0048: data <= 32'h133A9793;	14'h0049: data <= 32'h137E6E7B;	14'h004A: data <= 32'h13C23FC8;	14'h004B: data <= 32'h14060B67;	14'h004C: data <= 32'h1449D144;	14'h004D: data <= 32'h148D914D;	14'h004E: data <= 32'h14D14B6C;	14'h004F: data <= 32'h1514FF90;	14'h0050: data <= 32'h1558ADA4;	14'h0051: data <= 32'h159C5595;	14'h0052: data <= 32'h15DFF750;	14'h0053: data <= 32'h162392C1;	14'h0054: data <= 32'h166727D4;	14'h0055: data <= 32'h16AAB677;	14'h0056: data <= 32'h16EE3E96;	14'h0057: data <= 32'h1731C01E;	14'h0058: data <= 32'h17753AFA;	14'h0059: data <= 32'h17B8AF18;	14'h005A: data <= 32'h17FC1C64;	14'h005B: data <= 32'h183F82CC;	14'h005C: data <= 32'h1882E23A;	14'h005D: data <= 32'h18C63A9D;	14'h005E: data <= 32'h19098BE1;	14'h005F: data <= 32'h194CD5F2;	14'h0060: data <= 32'h199018BD;	14'h0061: data <= 32'h19D3542F;	14'h0062: data <= 32'h1A168834;	14'h0063: data <= 32'h1A59B4B9;	14'h0064: data <= 32'h1A9CD9AC;	14'h0065: data <= 32'h1ADFF6F7;	14'h0066: data <= 32'h1B230C89;	14'h0067: data <= 32'h1B661A4E;	14'h0068: data <= 32'h1BA92032;	14'h0069: data <= 32'h1BEC1E23;	14'h006A: data <= 32'h1C2F140D;	14'h006B: data <= 32'h1C7201DD;	14'h006C: data <= 32'h1CB4E77F;	14'h006D: data <= 32'h1CF7C4E1;	14'h006E: data <= 32'h1D3A99EF;	14'h006F: data <= 32'h1D7D6696;	14'h0070: data <= 32'h1DC02AC2;	14'h0071: data <= 32'h1E02E662;	14'h0072: data <= 32'h1E459960;	14'h0073: data <= 32'h1E8843AB;	14'h0074: data <= 32'h1ECAE52F;	14'h0075: data <= 32'h1F0D7DD8;	14'h0076: data <= 32'h1F500D95;	14'h0077: data <= 32'h1F929451;	14'h0078: data <= 32'h1FD511F9;	14'h0079: data <= 32'h2017867B;	14'h007A: data <= 32'h2059F1C3;	14'h007B: data <= 32'h209C53BF;	14'h007C: data <= 32'h20DEAC5A;	14'h007D: data <= 32'h2120FB82;	14'h007E: data <= 32'h21634125;	14'h007F: data <= 32'h21A57D2E;	14'h0080: data <= 32'h21E7AF8B;	14'h0081: data <= 32'h2229D829;	14'h0082: data <= 32'h226BF6F5;	14'h0083: data <= 32'h22AE0BDB;	14'h0084: data <= 32'h22F016C9;	14'h0085: data <= 32'h233217AD;	14'h0086: data <= 32'h23740E72;	14'h0087: data <= 32'h23B5FB05;	14'h0088: data <= 32'h23F7DD55;	14'h0089: data <= 32'h2439B54E;	14'h008A: data <= 32'h247B82DD;	14'h008B: data <= 32'h24BD45EF;	14'h008C: data <= 32'h24FEFE71;	14'h008D: data <= 32'h2540AC50;	14'h008E: data <= 32'h25824F7A;	14'h008F: data <= 32'h25C3E7DC;	14'h0090: data <= 32'h26057562;	14'h0091: data <= 32'h2646F7FB;	14'h0092: data <= 32'h26886F92;	14'h0093: data <= 32'h26C9DC16;	14'h0094: data <= 32'h270B3D72;	14'h0095: data <= 32'h274C9396;	14'h0096: data <= 32'h278DDE6E;	14'h0097: data <= 32'h27CF1DE6;	14'h0098: data <= 32'h281051ED;	14'h0099: data <= 32'h28517A6F;	14'h009A: data <= 32'h2892975B;	14'h009B: data <= 32'h28D3A89C;	14'h009C: data <= 32'h2914AE21;	14'h009D: data <= 32'h2955A7D7;	14'h009E: data <= 32'h299695AA;	14'h009F: data <= 32'h29D7778A;	14'h00A0: data <= 32'h2A184D61;	14'h00A1: data <= 32'h2A59171F;	14'h00A2: data <= 32'h2A99D4B1;	14'h00A3: data <= 32'h2ADA8603;	14'h00A4: data <= 32'h2B1B2B04;	14'h00A5: data <= 32'h2B5BC3A0;	14'h00A6: data <= 32'h2B9C4FC5;	14'h00A7: data <= 32'h2BDCCF61;	14'h00A8: data <= 32'h2C1D4261;	14'h00A9: data <= 32'h2C5DA8B3;	14'h00AA: data <= 32'h2C9E0243;	14'h00AB: data <= 32'h2CDE4F00;	14'h00AC: data <= 32'h2D1E8ED7;	14'h00AD: data <= 32'h2D5EC1B5;	14'h00AE: data <= 32'h2D9EE789;	14'h00AF: data <= 32'h2DDF003F;	14'h00B0: data <= 32'h2E1F0BC5;	14'h00B1: data <= 32'h2E5F0A09;	14'h00B2: data <= 32'h2E9EFAF9;	14'h00B3: data <= 32'h2EDEDE81;	14'h00B4: data <= 32'h2F1EB490;	14'h00B5: data <= 32'h2F5E7D14;	14'h00B6: data <= 32'h2F9E37F9;	14'h00B7: data <= 32'h2FDDE52E;	14'h00B8: data <= 32'h301D84A1;	14'h00B9: data <= 32'h305D163E;	14'h00BA: data <= 32'h309C99F5;	14'h00BB: data <= 32'h30DC0FB1;	14'h00BC: data <= 32'h311B7762;	14'h00BD: data <= 32'h315AD0F5;	14'h00BE: data <= 32'h319A1C58;	14'h00BF: data <= 32'h31D95979;	14'h00C0: data <= 32'h32188845;	14'h00C1: data <= 32'h3257A8AA;	14'h00C2: data <= 32'h3296BA97;	14'h00C3: data <= 32'h32D5BDF8;	14'h00C4: data <= 32'h3314B2BC;	14'h00C5: data <= 32'h335398D2;	14'h00C6: data <= 32'h33927025;	14'h00C7: data <= 32'h33D138A6;	14'h00C8: data <= 32'h340FF241;	14'h00C9: data <= 32'h344E9CE5;	14'h00CA: data <= 32'h348D387F;	14'h00CB: data <= 32'h34CBC4FE;	14'h00CC: data <= 32'h350A424F;	14'h00CD: data <= 32'h3548B061;	14'h00CE: data <= 32'h35870F22;	14'h00CF: data <= 32'h35C55E80;	14'h00D0: data <= 32'h36039E68;	14'h00D1: data <= 32'h3641CEC9;	14'h00D2: data <= 32'h367FEF91;	14'h00D3: data <= 32'h36BE00AF;	14'h00D4: data <= 32'h36FC0210;	14'h00D5: data <= 32'h3739F3A2;	14'h00D6: data <= 32'h3777D554;	14'h00D7: data <= 32'h37B5A714;	14'h00D8: data <= 32'h37F368D0;	14'h00D9: data <= 32'h38311A77;	14'h00DA: data <= 32'h386EBBF6;	14'h00DB: data <= 32'h38AC4D3C;	14'h00DC: data <= 32'h38E9CE38;	14'h00DD: data <= 32'h39273ED7;	14'h00DE: data <= 32'h39649F08;	14'h00DF: data <= 32'h39A1EEB9;	14'h00E0: data <= 32'h39DF2DD9;	14'h00E1: data <= 32'h3A1C5C56;	14'h00E2: data <= 32'h3A597A1E;	14'h00E3: data <= 32'h3A968720;	14'h00E4: data <= 32'h3AD3834B;	14'h00E5: data <= 32'h3B106E8C;	14'h00E6: data <= 32'h3B4D48D3;	14'h00E7: data <= 32'h3B8A120D;	14'h00E8: data <= 32'h3BC6CA2A;	14'h00E9: data <= 32'h3C037117;	14'h00EA: data <= 32'h3C4006C4;	14'h00EB: data <= 32'h3C7C8B1F;	14'h00EC: data <= 32'h3CB8FE17;	14'h00ED: data <= 32'h3CF55F9A;	14'h00EE: data <= 32'h3D31AF97;	14'h00EF: data <= 32'h3D6DEDFC;	14'h00F0: data <= 32'h3DAA1AB9;	14'h00F1: data <= 32'h3DE635BB;	14'h00F2: data <= 32'h3E223EF2;	14'h00F3: data <= 32'h3E5E364C;	14'h00F4: data <= 32'h3E9A1BB9;	14'h00F5: data <= 32'h3ED5EF27;	14'h00F6: data <= 32'h3F11B084;	14'h00F7: data <= 32'h3F4D5FC0;	14'h00F8: data <= 32'h3F88FCC9;	14'h00F9: data <= 32'h3FC4878E;	14'h00FA: data <= 32'h3FFFFFFF;	14'h00FB: data <= 32'h403B660A;	14'h00FC: data <= 32'h4076B99D;	14'h00FD: data <= 32'h40B1FAA9;	14'h00FE: data <= 32'h40ED291B;	14'h00FF: data <= 32'h412844E3;	14'h0100: data <= 32'h41634DF1;	14'h0101: data <= 32'h419E4432;	14'h0102: data <= 32'h41D92796;	14'h0103: data <= 32'h4213F80C;	14'h0104: data <= 32'h424EB583;	14'h0105: data <= 32'h42895FEA;	14'h0106: data <= 32'h42C3F731;	14'h0107: data <= 32'h42FE7B46;	14'h0108: data <= 32'h4338EC19;	14'h0109: data <= 32'h43734999;	14'h010A: data <= 32'h43AD93B5;	14'h010B: data <= 32'h43E7CA5C;	14'h010C: data <= 32'h4421ED7E;	14'h010D: data <= 32'h445BFD0A;	14'h010E: data <= 32'h4495F8EF;	14'h010F: data <= 32'h44CFE11D;	14'h0110: data <= 32'h4509B583;	14'h0111: data <= 32'h4543760F;	14'h0112: data <= 32'h457D22B3;	14'h0113: data <= 32'h45B6BB5D;	14'h0114: data <= 32'h45F03FFC;	14'h0115: data <= 32'h4629B080;	14'h0116: data <= 32'h46630CD9;	14'h0117: data <= 32'h469C54F6;	14'h0118: data <= 32'h46D588C6;	14'h0119: data <= 32'h470EA839;	14'h011A: data <= 32'h4747B33F;	14'h011B: data <= 32'h4780A9C8;	14'h011C: data <= 32'h47B98BC2;	14'h011D: data <= 32'h47F2591E;	14'h011E: data <= 32'h482B11CB;	14'h011F: data <= 32'h4863B5B9;	14'h0120: data <= 32'h489C44D7;	14'h0121: data <= 32'h48D4BF16;	14'h0122: data <= 32'h490D2465;	14'h0123: data <= 32'h494574B4;	14'h0124: data <= 32'h497DAFF3;	14'h0125: data <= 32'h49B5D611;	14'h0126: data <= 32'h49EDE6FF;	14'h0127: data <= 32'h4A25E2AC;	14'h0128: data <= 32'h4A5DC908;	14'h0129: data <= 32'h4A959A04;	14'h012A: data <= 32'h4ACD558E;	14'h012B: data <= 32'h4B04FB98;	14'h012C: data <= 32'h4B3C8C11;	14'h012D: data <= 32'h4B7406E9;	14'h012E: data <= 32'h4BAB6C10;	14'h012F: data <= 32'h4BE2BB76;	14'h0130: data <= 32'h4C19F50B;	14'h0131: data <= 32'h4C5118C0;	14'h0132: data <= 32'h4C882685;	14'h0133: data <= 32'h4CBF1E4A;	14'h0134: data <= 32'h4CF5FFFE;	14'h0135: data <= 32'h4D2CCB93;	14'h0136: data <= 32'h4D6380F8;	14'h0137: data <= 32'h4D9A201D;	14'h0138: data <= 32'h4DD0A8F4;	14'h0139: data <= 32'h4E071B6D;	14'h013A: data <= 32'h4E3D7776;	14'h013B: data <= 32'h4E73BD02;	14'h013C: data <= 32'h4EA9EC01;	14'h013D: data <= 32'h4EE00462;	14'h013E: data <= 32'h4F160617;	14'h013F: data <= 32'h4F4BF10F;	14'h0140: data <= 32'h4F81C53C;	14'h0141: data <= 32'h4FB7828E;	14'h0142: data <= 32'h4FED28F5;	14'h0143: data <= 32'h5022B862;	14'h0144: data <= 32'h505830C5;	14'h0145: data <= 32'h508D9210;	14'h0146: data <= 32'h50C2DC33;	14'h0147: data <= 32'h50F80F1E;	14'h0148: data <= 32'h512D2AC2;	14'h0149: data <= 32'h51622F11;	14'h014A: data <= 32'h51971BFA;	14'h014B: data <= 32'h51CBF16E;	14'h014C: data <= 32'h5200AF5F;	14'h014D: data <= 32'h523555BD;	14'h014E: data <= 32'h5269E47A;	14'h014F: data <= 32'h529E5B85;	14'h0150: data <= 32'h52D2BAD0;	14'h0151: data <= 32'h5307024B;	14'h0152: data <= 32'h533B31E9;	14'h0153: data <= 32'h536F4999;	14'h0154: data <= 32'h53A3494D;	14'h0155: data <= 32'h53D730F6;	14'h0156: data <= 32'h540B0085;	14'h0157: data <= 32'h543EB7EB;	14'h0158: data <= 32'h54725719;	14'h0159: data <= 32'h54A5DE00;	14'h015A: data <= 32'h54D94C92;	14'h015B: data <= 32'h550CA2BF;	14'h015C: data <= 32'h553FE07A;	14'h015D: data <= 32'h557305B2;	14'h015E: data <= 32'h55A6125A;	14'h015F: data <= 32'h55D90663;	14'h0160: data <= 32'h560BE1BF;	14'h0161: data <= 32'h563EA45D;	14'h0162: data <= 32'h56714E31;	14'h0163: data <= 32'h56A3DF2B;	14'h0164: data <= 32'h56D6573E;	14'h0165: data <= 32'h5708B659;	14'h0166: data <= 32'h573AFC6F;	14'h0167: data <= 32'h576D2972;	14'h0168: data <= 32'h579F3D53;	14'h0169: data <= 32'h57D13804;	14'h016A: data <= 32'h58031975;	14'h016B: data <= 32'h5834E19A;	14'h016C: data <= 32'h58669063;	14'h016D: data <= 32'h589825C3;	14'h016E: data <= 32'h58C9A1AA;	14'h016F: data <= 32'h58FB040C;	14'h0170: data <= 32'h592C4CD9;	14'h0171: data <= 32'h595D7C04;	14'h0172: data <= 32'h598E917E;	14'h0173: data <= 32'h59BF8D39;	14'h0174: data <= 32'h59F06F27;	14'h0175: data <= 32'h5A21373B;	14'h0176: data <= 32'h5A51E565;	14'h0177: data <= 32'h5A827999;	14'h0178: data <= 32'h5AB2F3C7;	14'h0179: data <= 32'h5AE353E3;	14'h017A: data <= 32'h5B1399DF;	14'h017B: data <= 32'h5B43C5AB;	14'h017C: data <= 32'h5B73D73B;	14'h017D: data <= 32'h5BA3CE81;	14'h017E: data <= 32'h5BD3AB6F;	14'h017F: data <= 32'h5C036DF7;	14'h0180: data <= 32'h5C33160B;	14'h0181: data <= 32'h5C62A39E;	14'h0182: data <= 32'h5C9216A3;	14'h0183: data <= 32'h5CC16F0A;	14'h0184: data <= 32'h5CF0ACC8;	14'h0185: data <= 32'h5D1FCFCE;	14'h0186: data <= 32'h5D4ED80E;	14'h0187: data <= 32'h5D7DC57C;	14'h0188: data <= 32'h5DAC9809;	14'h0189: data <= 32'h5DDB4FA9;	14'h018A: data <= 32'h5E09EC4D;	14'h018B: data <= 32'h5E386DE9;	14'h018C: data <= 32'h5E66D46E;	14'h018D: data <= 32'h5E951FD1;	14'h018E: data <= 32'h5EC35003;	14'h018F: data <= 32'h5EF164F7;	14'h0190: data <= 32'h5F1F5EA0;	14'h0191: data <= 32'h5F4D3CF0;	14'h0192: data <= 32'h5F7AFFDB;	14'h0193: data <= 32'h5FA8A753;	14'h0194: data <= 32'h5FD6334C;	14'h0195: data <= 32'h6003A3B7;	14'h0196: data <= 32'h6030F888;	14'h0197: data <= 32'h605E31B3;	14'h0198: data <= 32'h608B4F29;	14'h0199: data <= 32'h60B850DF;	14'h019A: data <= 32'h60E536C6;	14'h019B: data <= 32'h611200D3;	14'h019C: data <= 32'h613EAEF8;	14'h019D: data <= 32'h616B4129;	14'h019E: data <= 32'h6197B758;	14'h019F: data <= 32'h61C41179;	14'h01A0: data <= 32'h61F04F7F;	14'h01A1: data <= 32'h621C715D;	14'h01A2: data <= 32'h62487707;	14'h01A3: data <= 32'h62746071;	14'h01A4: data <= 32'h62A02D8C;	14'h01A5: data <= 32'h62CBDE4E;	14'h01A6: data <= 32'h62F772A8;	14'h01A7: data <= 32'h6322EA90;	14'h01A8: data <= 32'h634E45F8;	14'h01A9: data <= 32'h637984D3;	14'h01AA: data <= 32'h63A4A716;	14'h01AB: data <= 32'h63CFACB4;	14'h01AC: data <= 32'h63FA95A0;	14'h01AD: data <= 32'h642561CF;	14'h01AE: data <= 32'h64501133;	14'h01AF: data <= 32'h647AA3C2;	14'h01B0: data <= 32'h64A5196D;	14'h01B1: data <= 32'h64CF722A;	14'h01B2: data <= 32'h64F9ADEC;	14'h01B3: data <= 32'h6523CCA7;	14'h01B4: data <= 32'h654DCE4F;	14'h01B5: data <= 32'h6577B2D7;	14'h01B6: data <= 32'h65A17A34;	14'h01B7: data <= 32'h65CB245A;	14'h01B8: data <= 32'h65F4B13D;	14'h01B9: data <= 32'h661E20D0;	14'h01BA: data <= 32'h66477308;	14'h01BB: data <= 32'h6670A7D9;	14'h01BC: data <= 32'h6699BF37;	14'h01BD: data <= 32'h66C2B917;	14'h01BE: data <= 32'h66EB956C;	14'h01BF: data <= 32'h6714542B;	14'h01C0: data <= 32'h673CF548;	14'h01C1: data <= 32'h676578B7;	14'h01C2: data <= 32'h678DDE6D;	14'h01C3: data <= 32'h67B6265E;	14'h01C4: data <= 32'h67DE507F;	14'h01C5: data <= 32'h68065CC4;	14'h01C6: data <= 32'h682E4B21;	14'h01C7: data <= 32'h68561B8B;	14'h01C8: data <= 32'h687DCDF7;	14'h01C9: data <= 32'h68A56259;	14'h01CA: data <= 32'h68CCD8A5;	14'h01CB: data <= 32'h68F430D2;	14'h01CC: data <= 32'h691B6AD2;	14'h01CD: data <= 32'h6942869B;	14'h01CE: data <= 32'h69698422;	14'h01CF: data <= 32'h6990635B;	14'h01D0: data <= 32'h69B7243B;	14'h01D1: data <= 32'h69DDC6B8;	14'h01D2: data <= 32'h6A044AC5;	14'h01D3: data <= 32'h6A2AB058;	14'h01D4: data <= 32'h6A50F766;	14'h01D5: data <= 32'h6A771FE4;	14'h01D6: data <= 32'h6A9D29C7;	14'h01D7: data <= 32'h6AC31504;	14'h01D8: data <= 32'h6AE8E190;	14'h01D9: data <= 32'h6B0E8F60;	14'h01DA: data <= 32'h6B341E69;	14'h01DB: data <= 32'h6B598EA1;	14'h01DC: data <= 32'h6B7EDFFD;	14'h01DD: data <= 32'h6BA41272;	14'h01DE: data <= 32'h6BC925F5;	14'h01DF: data <= 32'h6BEE1A7C;	14'h01E0: data <= 32'h6C12EFFC;	14'h01E1: data <= 32'h6C37A66B;	14'h01E2: data <= 32'h6C5C3DBD;	14'h01E3: data <= 32'h6C80B5E9;	14'h01E4: data <= 32'h6CA50EE4;	14'h01E5: data <= 32'h6CC948A3;	14'h01E6: data <= 32'h6CED631D;	14'h01E7: data <= 32'h6D115E46;	14'h01E8: data <= 32'h6D353A15;	14'h01E9: data <= 32'h6D58F67E;	14'h01EA: data <= 32'h6D7C9378;	14'h01EB: data <= 32'h6DA010F9;	14'h01EC: data <= 32'h6DC36EF7;	14'h01ED: data <= 32'h6DE6AD66;	14'h01EE: data <= 32'h6E09CC3D;	14'h01EF: data <= 32'h6E2CCB73;	14'h01F0: data <= 32'h6E4FAAFC;	14'h01F1: data <= 32'h6E726ACF;	14'h01F2: data <= 32'h6E950AE2;	14'h01F3: data <= 32'h6EB78B2B;	14'h01F4: data <= 32'h6ED9EBA0;	14'h01F5: data <= 32'h6EFC2C37;	14'h01F6: data <= 32'h6F1E4CE6;	14'h01F7: data <= 32'h6F404DA4;	14'h01F8: data <= 32'h6F622E67;	14'h01F9: data <= 32'h6F83EF24;	14'h01FA: data <= 32'h6FA58FD3;	14'h01FB: data <= 32'h6FC71069;	14'h01FC: data <= 32'h6FE870DD;	14'h01FD: data <= 32'h7009B125;	14'h01FE: data <= 32'h702AD139;	14'h01FF: data <= 32'h704BD10D;	14'h0200: data <= 32'h706CB09A;	14'h0201: data <= 32'h708D6FD4;	14'h0202: data <= 32'h70AE0EB4;	14'h0203: data <= 32'h70CE8D2F;	14'h0204: data <= 32'h70EEEB3C;	14'h0205: data <= 32'h710F28D2;	14'h0206: data <= 32'h712F45E8;	14'h0207: data <= 32'h714F4274;	14'h0208: data <= 32'h716F1E6E;	14'h0209: data <= 32'h718ED9CB;	14'h020A: data <= 32'h71AE7484;	14'h020B: data <= 32'h71CDEE8E;	14'h020C: data <= 32'h71ED47E1;	14'h020D: data <= 32'h720C8074;	14'h020E: data <= 32'h722B983D;	14'h020F: data <= 32'h724A8F35;	14'h0210: data <= 32'h72696551;	14'h0211: data <= 32'h72881A89;	14'h0212: data <= 32'h72A6AED5;	14'h0213: data <= 32'h72C5222B;	14'h0214: data <= 32'h72E37483;	14'h0215: data <= 32'h7301A5D4;	14'h0216: data <= 32'h731FB615;	14'h0217: data <= 32'h733DA53E;	14'h0218: data <= 32'h735B7346;	14'h0219: data <= 32'h73792025;	14'h021A: data <= 32'h7396ABD1;	14'h021B: data <= 32'h73B41643;	14'h021C: data <= 32'h73D15F72;	14'h021D: data <= 32'h73EE8756;	14'h021E: data <= 32'h740B8DE5;	14'h021F: data <= 32'h74287319;	14'h0220: data <= 32'h744536E8;	14'h0221: data <= 32'h7461D94B;	14'h0222: data <= 32'h747E5A39;	14'h0223: data <= 32'h749AB9A9;	14'h0224: data <= 32'h74B6F794;	14'h0225: data <= 32'h74D313F2;	14'h0226: data <= 32'h74EF0EBB;	14'h0227: data <= 32'h750AE7E5;	14'h0228: data <= 32'h75269F6B;	14'h0229: data <= 32'h75423543;	14'h022A: data <= 32'h755DA965;	14'h022B: data <= 32'h7578FBCA;	14'h022C: data <= 32'h75942C6A;	14'h022D: data <= 32'h75AF3B3D;	14'h022E: data <= 32'h75CA283B;	14'h022F: data <= 32'h75E4F35D;	14'h0230: data <= 32'h75FF9C9A;	14'h0231: data <= 32'h761A23EC;	14'h0232: data <= 32'h7634894A;	14'h0233: data <= 32'h764ECCAD;	14'h0234: data <= 32'h7668EE0D;	14'h0235: data <= 32'h7682ED64;	14'h0236: data <= 32'h769CCAA8;	14'h0237: data <= 32'h76B685D4;	14'h0238: data <= 32'h76D01EDF;	14'h0239: data <= 32'h76E995C2;	14'h023A: data <= 32'h7702EA76;	14'h023B: data <= 32'h771C1CF4;	14'h023C: data <= 32'h77352D34;	14'h023D: data <= 32'h774E1B2F;	14'h023E: data <= 32'h7766E6DF;	14'h023F: data <= 32'h777F903B;	14'h0240: data <= 32'h7798173C;	14'h0241: data <= 32'h77B07BDD;	14'h0242: data <= 32'h77C8BE15;	14'h0243: data <= 32'h77E0DDDE;	14'h0244: data <= 32'h77F8DB31;	14'h0245: data <= 32'h7810B606;	14'h0246: data <= 32'h78286E58;	14'h0247: data <= 32'h7840041E;	14'h0248: data <= 32'h78577754;	14'h0249: data <= 32'h786EC7F1;	14'h024A: data <= 32'h7885F5EE;	14'h024B: data <= 32'h789D0147;	14'h024C: data <= 32'h78B3E9F3;	14'h024D: data <= 32'h78CAAFEC;	14'h024E: data <= 32'h78E1532B;	14'h024F: data <= 32'h78F7D3AB;	14'h0250: data <= 32'h790E3164;	14'h0251: data <= 32'h79246C50;	14'h0252: data <= 32'h793A846A;	14'h0253: data <= 32'h795079A9;	14'h0254: data <= 32'h79664C09;	14'h0255: data <= 32'h797BFB82;	14'h0256: data <= 32'h7991880F;	14'h0257: data <= 32'h79A6F1AA;	14'h0258: data <= 32'h79BC384C;	14'h0259: data <= 32'h79D15BEE;	14'h025A: data <= 32'h79E65C8C;	14'h025B: data <= 32'h79FB3A1F;	14'h025C: data <= 32'h7A0FF4A1;	14'h025D: data <= 32'h7A248C0C;	14'h025E: data <= 32'h7A39005A;	14'h025F: data <= 32'h7A4D5186;	14'h0260: data <= 32'h7A617F89;	14'h0261: data <= 32'h7A758A5D;	14'h0262: data <= 32'h7A8971FD;	14'h0263: data <= 32'h7A9D3664;	14'h0264: data <= 32'h7AB0D78B;	14'h0265: data <= 32'h7AC4556C;	14'h0266: data <= 32'h7AD7B003;	14'h0267: data <= 32'h7AEAE74A;	14'h0268: data <= 32'h7AFDFB3A;	14'h0269: data <= 32'h7B10EBD0;	14'h026A: data <= 32'h7B23B904;	14'h026B: data <= 32'h7B3662D2;	14'h026C: data <= 32'h7B48E935;	14'h026D: data <= 32'h7B5B4C27;	14'h026E: data <= 32'h7B6D8BA2;	14'h026F: data <= 32'h7B7FA7A3;	14'h0270: data <= 32'h7B91A022;	14'h0271: data <= 32'h7BA3751C;	14'h0272: data <= 32'h7BB5268A;	14'h0273: data <= 32'h7BC6B469;	14'h0274: data <= 32'h7BD81EB3;	14'h0275: data <= 32'h7BE96562;	14'h0276: data <= 32'h7BFA8873;	14'h0277: data <= 32'h7C0B87DF;	14'h0278: data <= 32'h7C1C63A3;	14'h0279: data <= 32'h7C2D1BB9;	14'h027A: data <= 32'h7C3DB01C;	14'h027B: data <= 32'h7C4E20C9;	14'h027C: data <= 32'h7C5E6DB9;	14'h027D: data <= 32'h7C6E96E8;	14'h027E: data <= 32'h7C7E9C53;	14'h027F: data <= 32'h7C8E7DF3;	14'h0280: data <= 32'h7C9E3BC4;	14'h0281: data <= 32'h7CADD5C3;	14'h0282: data <= 32'h7CBD4BEA;	14'h0283: data <= 32'h7CCC9E36;	14'h0284: data <= 32'h7CDBCCA0;	14'h0285: data <= 32'h7CEAD727;	14'h0286: data <= 32'h7CF9BDC4;	14'h0287: data <= 32'h7D088073;	14'h0288: data <= 32'h7D171F32;	14'h0289: data <= 32'h7D2599FA;	14'h028A: data <= 32'h7D33F0C8;	14'h028B: data <= 32'h7D422399;	14'h028C: data <= 32'h7D503267;	14'h028D: data <= 32'h7D5E1D2F;	14'h028E: data <= 32'h7D6BE3ED;	14'h028F: data <= 32'h7D79869D;	14'h0290: data <= 32'h7D87053A;	14'h0291: data <= 32'h7D945FC2;	14'h0292: data <= 32'h7DA19630;	14'h0293: data <= 32'h7DAEA880;	14'h0294: data <= 32'h7DBB96AF;	14'h0295: data <= 32'h7DC860B9;	14'h0296: data <= 32'h7DD5069A;	14'h0297: data <= 32'h7DE1884F;	14'h0298: data <= 32'h7DEDE5D4;	14'h0299: data <= 32'h7DFA1F25;	14'h029A: data <= 32'h7E06343F;	14'h029B: data <= 32'h7E12251F;	14'h029C: data <= 32'h7E1DF1C1;	14'h029D: data <= 32'h7E299A21;	14'h029E: data <= 32'h7E351E3D;	14'h029F: data <= 32'h7E407E11;	14'h02A0: data <= 32'h7E4BB999;	14'h02A1: data <= 32'h7E56D0D3;	14'h02A2: data <= 32'h7E61C3BC;	14'h02A3: data <= 32'h7E6C924F;	14'h02A4: data <= 32'h7E773C8B;	14'h02A5: data <= 32'h7E81C26B;	14'h02A6: data <= 32'h7E8C23EE;	14'h02A7: data <= 32'h7E96610F;	14'h02A8: data <= 32'h7EA079CD;	14'h02A9: data <= 32'h7EAA6E24;	14'h02AA: data <= 32'h7EB43E11;	14'h02AB: data <= 32'h7EBDE991;	14'h02AC: data <= 32'h7EC770A2;	14'h02AD: data <= 32'h7ED0D341;	14'h02AE: data <= 32'h7EDA116B;	14'h02AF: data <= 32'h7EE32B1E;	14'h02B0: data <= 32'h7EEC2057;	14'h02B1: data <= 32'h7EF4F113;	14'h02B2: data <= 32'h7EFD9D51;	14'h02B3: data <= 32'h7F06250C;	14'h02B4: data <= 32'h7F0E8843;	14'h02B5: data <= 32'h7F16C6F4;	14'h02B6: data <= 32'h7F1EE11C;	14'h02B7: data <= 32'h7F26D6B9;	14'h02B8: data <= 32'h7F2EA7C8;	14'h02B9: data <= 32'h7F365448;	14'h02BA: data <= 32'h7F3DDC36;	14'h02BB: data <= 32'h7F453F8F;	14'h02BC: data <= 32'h7F4C7E52;	14'h02BD: data <= 32'h7F53987D;	14'h02BE: data <= 32'h7F5A8E0E;	14'h02BF: data <= 32'h7F615F02;	14'h02C0: data <= 32'h7F680B58;	14'h02C1: data <= 32'h7F6E930E;	14'h02C2: data <= 32'h7F74F622;	14'h02C3: data <= 32'h7F7B3491;	14'h02C4: data <= 32'h7F814E5B;	14'h02C5: data <= 32'h7F87437E;	14'h02C6: data <= 32'h7F8D13F7;	14'h02C7: data <= 32'h7F92BFC5;	14'h02C8: data <= 32'h7F9846E7;	14'h02C9: data <= 32'h7F9DA95B;	14'h02CA: data <= 32'h7FA2E71F;	14'h02CB: data <= 32'h7FA80032;	14'h02CC: data <= 32'h7FACF493;	14'h02CD: data <= 32'h7FB1C43F;	14'h02CE: data <= 32'h7FB66F36;	14'h02CF: data <= 32'h7FBAF576;	14'h02D0: data <= 32'h7FBF56FE;	14'h02D1: data <= 32'h7FC393CD;	14'h02D2: data <= 32'h7FC7ABE1;	14'h02D3: data <= 32'h7FCB9F39;	14'h02D4: data <= 32'h7FCF6DD5;	14'h02D5: data <= 32'h7FD317B3;	14'h02D6: data <= 32'h7FD69CD1;	14'h02D7: data <= 32'h7FD9FD30;	14'h02D8: data <= 32'h7FDD38CE;	14'h02D9: data <= 32'h7FE04FAA;	14'h02DA: data <= 32'h7FE341C2;	14'h02DB: data <= 32'h7FE60F18;	14'h02DC: data <= 32'h7FE8B7A9;	14'h02DD: data <= 32'h7FEB3B74;	14'h02DE: data <= 32'h7FED9A7A;	14'h02DF: data <= 32'h7FEFD4B9;	14'h02E0: data <= 32'h7FF1EA31;	14'h02E1: data <= 32'h7FF3DAE1;	14'h02E2: data <= 32'h7FF5A6C8;	14'h02E3: data <= 32'h7FF74DE7;	14'h02E4: data <= 32'h7FF8D03C;	14'h02E5: data <= 32'h7FFA2DC7;	14'h02E6: data <= 32'h7FFB6688;	14'h02E7: data <= 32'h7FFC7A7F;	14'h02E8: data <= 32'h7FFD69AA;	14'h02E9: data <= 32'h7FFE340B;	14'h02EA: data <= 32'h7FFED9A0;	14'h02EB: data <= 32'h7FFF5A69;	14'h02EC: data <= 32'h7FFFB667;	14'h02ED: data <= 32'h7FFFED99;	14'h02EE: data <= 32'h7FFFFFFF;	14'h02EF: data <= 32'h7FFFED99;	14'h02F0: data <= 32'h7FFFB667;	14'h02F1: data <= 32'h7FFF5A69;	14'h02F2: data <= 32'h7FFED9A0;	14'h02F3: data <= 32'h7FFE340B;	14'h02F4: data <= 32'h7FFD69AA;	14'h02F5: data <= 32'h7FFC7A7F;	14'h02F6: data <= 32'h7FFB6688;	14'h02F7: data <= 32'h7FFA2DC7;	14'h02F8: data <= 32'h7FF8D03C;	14'h02F9: data <= 32'h7FF74DE7;	14'h02FA: data <= 32'h7FF5A6C8;	14'h02FB: data <= 32'h7FF3DAE1;	14'h02FC: data <= 32'h7FF1EA31;	14'h02FD: data <= 32'h7FEFD4B9;	14'h02FE: data <= 32'h7FED9A7A;	14'h02FF: data <= 32'h7FEB3B74;	14'h0300: data <= 32'h7FE8B7A9;	14'h0301: data <= 32'h7FE60F18;	14'h0302: data <= 32'h7FE341C2;	14'h0303: data <= 32'h7FE04FAA;	14'h0304: data <= 32'h7FDD38CE;	14'h0305: data <= 32'h7FD9FD30;	14'h0306: data <= 32'h7FD69CD1;	14'h0307: data <= 32'h7FD317B3;	14'h0308: data <= 32'h7FCF6DD5;	14'h0309: data <= 32'h7FCB9F39;	14'h030A: data <= 32'h7FC7ABE1;	14'h030B: data <= 32'h7FC393CD;	14'h030C: data <= 32'h7FBF56FE;	14'h030D: data <= 32'h7FBAF576;	14'h030E: data <= 32'h7FB66F36;	14'h030F: data <= 32'h7FB1C43F;	14'h0310: data <= 32'h7FACF493;	14'h0311: data <= 32'h7FA80032;	14'h0312: data <= 32'h7FA2E71F;	14'h0313: data <= 32'h7F9DA95B;	14'h0314: data <= 32'h7F9846E7;	14'h0315: data <= 32'h7F92BFC5;	14'h0316: data <= 32'h7F8D13F7;	14'h0317: data <= 32'h7F87437E;	14'h0318: data <= 32'h7F814E5B;	14'h0319: data <= 32'h7F7B3491;	14'h031A: data <= 32'h7F74F622;	14'h031B: data <= 32'h7F6E930E;	14'h031C: data <= 32'h7F680B58;	14'h031D: data <= 32'h7F615F02;	14'h031E: data <= 32'h7F5A8E0E;	14'h031F: data <= 32'h7F53987D;	14'h0320: data <= 32'h7F4C7E52;	14'h0321: data <= 32'h7F453F8F;	14'h0322: data <= 32'h7F3DDC36;	14'h0323: data <= 32'h7F365448;	14'h0324: data <= 32'h7F2EA7C8;	14'h0325: data <= 32'h7F26D6B9;	14'h0326: data <= 32'h7F1EE11C;	14'h0327: data <= 32'h7F16C6F4;	14'h0328: data <= 32'h7F0E8843;	14'h0329: data <= 32'h7F06250C;	14'h032A: data <= 32'h7EFD9D51;	14'h032B: data <= 32'h7EF4F113;	14'h032C: data <= 32'h7EEC2057;	14'h032D: data <= 32'h7EE32B1E;	14'h032E: data <= 32'h7EDA116B;	14'h032F: data <= 32'h7ED0D341;	14'h0330: data <= 32'h7EC770A2;	14'h0331: data <= 32'h7EBDE991;	14'h0332: data <= 32'h7EB43E11;	14'h0333: data <= 32'h7EAA6E24;	14'h0334: data <= 32'h7EA079CD;	14'h0335: data <= 32'h7E96610F;	14'h0336: data <= 32'h7E8C23EE;	14'h0337: data <= 32'h7E81C26B;	14'h0338: data <= 32'h7E773C8B;	14'h0339: data <= 32'h7E6C924F;	14'h033A: data <= 32'h7E61C3BC;	14'h033B: data <= 32'h7E56D0D3;	14'h033C: data <= 32'h7E4BB999;	14'h033D: data <= 32'h7E407E11;	14'h033E: data <= 32'h7E351E3D;	14'h033F: data <= 32'h7E299A21;	14'h0340: data <= 32'h7E1DF1C1;	14'h0341: data <= 32'h7E12251F;	14'h0342: data <= 32'h7E06343F;	14'h0343: data <= 32'h7DFA1F25;	14'h0344: data <= 32'h7DEDE5D4;	14'h0345: data <= 32'h7DE1884F;	14'h0346: data <= 32'h7DD5069A;	14'h0347: data <= 32'h7DC860B9;	14'h0348: data <= 32'h7DBB96AF;	14'h0349: data <= 32'h7DAEA880;	14'h034A: data <= 32'h7DA19630;	14'h034B: data <= 32'h7D945FC2;	14'h034C: data <= 32'h7D87053A;	14'h034D: data <= 32'h7D79869D;	14'h034E: data <= 32'h7D6BE3ED;	14'h034F: data <= 32'h7D5E1D2F;	14'h0350: data <= 32'h7D503267;	14'h0351: data <= 32'h7D422399;	14'h0352: data <= 32'h7D33F0C8;	14'h0353: data <= 32'h7D2599FA;	14'h0354: data <= 32'h7D171F32;	14'h0355: data <= 32'h7D088073;	14'h0356: data <= 32'h7CF9BDC4;	14'h0357: data <= 32'h7CEAD727;	14'h0358: data <= 32'h7CDBCCA0;	14'h0359: data <= 32'h7CCC9E36;	14'h035A: data <= 32'h7CBD4BEA;	14'h035B: data <= 32'h7CADD5C3;	14'h035C: data <= 32'h7C9E3BC4;	14'h035D: data <= 32'h7C8E7DF3;	14'h035E: data <= 32'h7C7E9C53;	14'h035F: data <= 32'h7C6E96E8;	14'h0360: data <= 32'h7C5E6DB9;	14'h0361: data <= 32'h7C4E20C9;	14'h0362: data <= 32'h7C3DB01C;	14'h0363: data <= 32'h7C2D1BB9;	14'h0364: data <= 32'h7C1C63A3;	14'h0365: data <= 32'h7C0B87DF;	14'h0366: data <= 32'h7BFA8873;	14'h0367: data <= 32'h7BE96562;	14'h0368: data <= 32'h7BD81EB3;	14'h0369: data <= 32'h7BC6B469;	14'h036A: data <= 32'h7BB5268A;	14'h036B: data <= 32'h7BA3751C;	14'h036C: data <= 32'h7B91A022;	14'h036D: data <= 32'h7B7FA7A3;	14'h036E: data <= 32'h7B6D8BA2;	14'h036F: data <= 32'h7B5B4C27;	14'h0370: data <= 32'h7B48E935;	14'h0371: data <= 32'h7B3662D2;	14'h0372: data <= 32'h7B23B904;	14'h0373: data <= 32'h7B10EBD0;	14'h0374: data <= 32'h7AFDFB3A;	14'h0375: data <= 32'h7AEAE74A;	14'h0376: data <= 32'h7AD7B003;	14'h0377: data <= 32'h7AC4556C;	14'h0378: data <= 32'h7AB0D78B;	14'h0379: data <= 32'h7A9D3664;	14'h037A: data <= 32'h7A8971FD;	14'h037B: data <= 32'h7A758A5D;	14'h037C: data <= 32'h7A617F89;	14'h037D: data <= 32'h7A4D5186;	14'h037E: data <= 32'h7A39005A;	14'h037F: data <= 32'h7A248C0C;	14'h0380: data <= 32'h7A0FF4A1;	14'h0381: data <= 32'h79FB3A1F;	14'h0382: data <= 32'h79E65C8C;	14'h0383: data <= 32'h79D15BEE;	14'h0384: data <= 32'h79BC384C;	14'h0385: data <= 32'h79A6F1AA;	14'h0386: data <= 32'h7991880F;	14'h0387: data <= 32'h797BFB82;	14'h0388: data <= 32'h79664C09;	14'h0389: data <= 32'h795079A9;	14'h038A: data <= 32'h793A846A;	14'h038B: data <= 32'h79246C50;	14'h038C: data <= 32'h790E3164;	14'h038D: data <= 32'h78F7D3AB;	14'h038E: data <= 32'h78E1532B;	14'h038F: data <= 32'h78CAAFEC;	14'h0390: data <= 32'h78B3E9F3;	14'h0391: data <= 32'h789D0147;	14'h0392: data <= 32'h7885F5EE;	14'h0393: data <= 32'h786EC7F1;	14'h0394: data <= 32'h78577754;	14'h0395: data <= 32'h7840041E;	14'h0396: data <= 32'h78286E58;	14'h0397: data <= 32'h7810B606;	14'h0398: data <= 32'h77F8DB31;	14'h0399: data <= 32'h77E0DDDE;	14'h039A: data <= 32'h77C8BE15;	14'h039B: data <= 32'h77B07BDD;	14'h039C: data <= 32'h7798173C;	14'h039D: data <= 32'h777F903B;	14'h039E: data <= 32'h7766E6DF;	14'h039F: data <= 32'h774E1B2F;	14'h03A0: data <= 32'h77352D34;	14'h03A1: data <= 32'h771C1CF4;	14'h03A2: data <= 32'h7702EA76;	14'h03A3: data <= 32'h76E995C2;	14'h03A4: data <= 32'h76D01EDF;	14'h03A5: data <= 32'h76B685D4;	14'h03A6: data <= 32'h769CCAA8;	14'h03A7: data <= 32'h7682ED64;	14'h03A8: data <= 32'h7668EE0D;	14'h03A9: data <= 32'h764ECCAD;	14'h03AA: data <= 32'h7634894A;	14'h03AB: data <= 32'h761A23EC;	14'h03AC: data <= 32'h75FF9C9A;	14'h03AD: data <= 32'h75E4F35D;	14'h03AE: data <= 32'h75CA283B;	14'h03AF: data <= 32'h75AF3B3D;	14'h03B0: data <= 32'h75942C6A;	14'h03B1: data <= 32'h7578FBCA;	14'h03B2: data <= 32'h755DA965;	14'h03B3: data <= 32'h75423543;	14'h03B4: data <= 32'h75269F6B;	14'h03B5: data <= 32'h750AE7E5;	14'h03B6: data <= 32'h74EF0EBB;	14'h03B7: data <= 32'h74D313F2;	14'h03B8: data <= 32'h74B6F794;	14'h03B9: data <= 32'h749AB9A9;	14'h03BA: data <= 32'h747E5A39;	14'h03BB: data <= 32'h7461D94B;	14'h03BC: data <= 32'h744536E8;	14'h03BD: data <= 32'h74287319;	14'h03BE: data <= 32'h740B8DE5;	14'h03BF: data <= 32'h73EE8756;	14'h03C0: data <= 32'h73D15F72;	14'h03C1: data <= 32'h73B41643;	14'h03C2: data <= 32'h7396ABD1;	14'h03C3: data <= 32'h73792025;	14'h03C4: data <= 32'h735B7346;	14'h03C5: data <= 32'h733DA53E;	14'h03C6: data <= 32'h731FB615;	14'h03C7: data <= 32'h7301A5D4;	14'h03C8: data <= 32'h72E37483;	14'h03C9: data <= 32'h72C5222B;	14'h03CA: data <= 32'h72A6AED5;	14'h03CB: data <= 32'h72881A89;	14'h03CC: data <= 32'h72696551;	14'h03CD: data <= 32'h724A8F35;	14'h03CE: data <= 32'h722B983D;	14'h03CF: data <= 32'h720C8074;	14'h03D0: data <= 32'h71ED47E1;	14'h03D1: data <= 32'h71CDEE8E;	14'h03D2: data <= 32'h71AE7484;	14'h03D3: data <= 32'h718ED9CB;	14'h03D4: data <= 32'h716F1E6E;	14'h03D5: data <= 32'h714F4274;	14'h03D6: data <= 32'h712F45E8;	14'h03D7: data <= 32'h710F28D2;	14'h03D8: data <= 32'h70EEEB3C;	14'h03D9: data <= 32'h70CE8D2F;	14'h03DA: data <= 32'h70AE0EB4;	14'h03DB: data <= 32'h708D6FD4;	14'h03DC: data <= 32'h706CB09A;	14'h03DD: data <= 32'h704BD10D;	14'h03DE: data <= 32'h702AD139;	14'h03DF: data <= 32'h7009B125;	14'h03E0: data <= 32'h6FE870DD;	14'h03E1: data <= 32'h6FC71069;	14'h03E2: data <= 32'h6FA58FD3;	14'h03E3: data <= 32'h6F83EF24;	14'h03E4: data <= 32'h6F622E67;	14'h03E5: data <= 32'h6F404DA4;	14'h03E6: data <= 32'h6F1E4CE6;	14'h03E7: data <= 32'h6EFC2C37;	14'h03E8: data <= 32'h6ED9EBA0;	14'h03E9: data <= 32'h6EB78B2B;	14'h03EA: data <= 32'h6E950AE2;	14'h03EB: data <= 32'h6E726ACF;	14'h03EC: data <= 32'h6E4FAAFC;	14'h03ED: data <= 32'h6E2CCB73;	14'h03EE: data <= 32'h6E09CC3D;	14'h03EF: data <= 32'h6DE6AD66;	14'h03F0: data <= 32'h6DC36EF7;	14'h03F1: data <= 32'h6DA010F9;	14'h03F2: data <= 32'h6D7C9378;	14'h03F3: data <= 32'h6D58F67E;	14'h03F4: data <= 32'h6D353A15;	14'h03F5: data <= 32'h6D115E46;	14'h03F6: data <= 32'h6CED631D;	14'h03F7: data <= 32'h6CC948A3;	14'h03F8: data <= 32'h6CA50EE4;	14'h03F9: data <= 32'h6C80B5E9;	14'h03FA: data <= 32'h6C5C3DBD;	14'h03FB: data <= 32'h6C37A66B;	14'h03FC: data <= 32'h6C12EFFC;	14'h03FD: data <= 32'h6BEE1A7C;	14'h03FE: data <= 32'h6BC925F5;	14'h03FF: data <= 32'h6BA41272;	14'h0400: data <= 32'h6B7EDFFD;	14'h0401: data <= 32'h6B598EA1;	14'h0402: data <= 32'h6B341E69;	14'h0403: data <= 32'h6B0E8F60;	14'h0404: data <= 32'h6AE8E190;	14'h0405: data <= 32'h6AC31504;	14'h0406: data <= 32'h6A9D29C7;	14'h0407: data <= 32'h6A771FE4;	14'h0408: data <= 32'h6A50F766;	14'h0409: data <= 32'h6A2AB058;	14'h040A: data <= 32'h6A044AC5;	14'h040B: data <= 32'h69DDC6B8;	14'h040C: data <= 32'h69B7243B;	14'h040D: data <= 32'h6990635B;	14'h040E: data <= 32'h69698422;	14'h040F: data <= 32'h6942869B;	14'h0410: data <= 32'h691B6AD2;	14'h0411: data <= 32'h68F430D2;	14'h0412: data <= 32'h68CCD8A5;	14'h0413: data <= 32'h68A56259;	14'h0414: data <= 32'h687DCDF7;	14'h0415: data <= 32'h68561B8B;	14'h0416: data <= 32'h682E4B21;	14'h0417: data <= 32'h68065CC4;	14'h0418: data <= 32'h67DE507F;	14'h0419: data <= 32'h67B6265E;	14'h041A: data <= 32'h678DDE6D;	14'h041B: data <= 32'h676578B7;	14'h041C: data <= 32'h673CF548;	14'h041D: data <= 32'h6714542B;	14'h041E: data <= 32'h66EB956C;	14'h041F: data <= 32'h66C2B917;	14'h0420: data <= 32'h6699BF37;	14'h0421: data <= 32'h6670A7D9;	14'h0422: data <= 32'h66477308;	14'h0423: data <= 32'h661E20D0;	14'h0424: data <= 32'h65F4B13D;	14'h0425: data <= 32'h65CB245A;	14'h0426: data <= 32'h65A17A34;	14'h0427: data <= 32'h6577B2D7;	14'h0428: data <= 32'h654DCE4F;	14'h0429: data <= 32'h6523CCA7;	14'h042A: data <= 32'h64F9ADEC;	14'h042B: data <= 32'h64CF722A;	14'h042C: data <= 32'h64A5196D;	14'h042D: data <= 32'h647AA3C2;	14'h042E: data <= 32'h64501133;	14'h042F: data <= 32'h642561CF;	14'h0430: data <= 32'h63FA95A0;	14'h0431: data <= 32'h63CFACB4;	14'h0432: data <= 32'h63A4A716;	14'h0433: data <= 32'h637984D3;	14'h0434: data <= 32'h634E45F8;	14'h0435: data <= 32'h6322EA90;	14'h0436: data <= 32'h62F772A8;	14'h0437: data <= 32'h62CBDE4E;	14'h0438: data <= 32'h62A02D8C;	14'h0439: data <= 32'h62746071;	14'h043A: data <= 32'h62487707;	14'h043B: data <= 32'h621C715D;	14'h043C: data <= 32'h61F04F7F;	14'h043D: data <= 32'h61C41179;	14'h043E: data <= 32'h6197B758;	14'h043F: data <= 32'h616B4129;	14'h0440: data <= 32'h613EAEF8;	14'h0441: data <= 32'h611200D3;	14'h0442: data <= 32'h60E536C6;	14'h0443: data <= 32'h60B850DF;	14'h0444: data <= 32'h608B4F29;	14'h0445: data <= 32'h605E31B3;	14'h0446: data <= 32'h6030F888;	14'h0447: data <= 32'h6003A3B7;	14'h0448: data <= 32'h5FD6334C;	14'h0449: data <= 32'h5FA8A753;	14'h044A: data <= 32'h5F7AFFDB;	14'h044B: data <= 32'h5F4D3CF0;	14'h044C: data <= 32'h5F1F5EA0;	14'h044D: data <= 32'h5EF164F7;	14'h044E: data <= 32'h5EC35003;	14'h044F: data <= 32'h5E951FD1;	14'h0450: data <= 32'h5E66D46E;	14'h0451: data <= 32'h5E386DE9;	14'h0452: data <= 32'h5E09EC4D;	14'h0453: data <= 32'h5DDB4FA9;	14'h0454: data <= 32'h5DAC9809;	14'h0455: data <= 32'h5D7DC57C;	14'h0456: data <= 32'h5D4ED80E;	14'h0457: data <= 32'h5D1FCFCE;	14'h0458: data <= 32'h5CF0ACC8;	14'h0459: data <= 32'h5CC16F0A;	14'h045A: data <= 32'h5C9216A3;	14'h045B: data <= 32'h5C62A39E;	14'h045C: data <= 32'h5C33160B;	14'h045D: data <= 32'h5C036DF7;	14'h045E: data <= 32'h5BD3AB6F;	14'h045F: data <= 32'h5BA3CE81;	14'h0460: data <= 32'h5B73D73B;	14'h0461: data <= 32'h5B43C5AB;	14'h0462: data <= 32'h5B1399DF;	14'h0463: data <= 32'h5AE353E3;	14'h0464: data <= 32'h5AB2F3C7;	14'h0465: data <= 32'h5A827999;	14'h0466: data <= 32'h5A51E565;	14'h0467: data <= 32'h5A21373B;	14'h0468: data <= 32'h59F06F27;	14'h0469: data <= 32'h59BF8D39;	14'h046A: data <= 32'h598E917E;	14'h046B: data <= 32'h595D7C04;	14'h046C: data <= 32'h592C4CD9;	14'h046D: data <= 32'h58FB040C;	14'h046E: data <= 32'h58C9A1AA;	14'h046F: data <= 32'h589825C3;	14'h0470: data <= 32'h58669063;	14'h0471: data <= 32'h5834E19A;	14'h0472: data <= 32'h58031975;	14'h0473: data <= 32'h57D13804;	14'h0474: data <= 32'h579F3D53;	14'h0475: data <= 32'h576D2972;	14'h0476: data <= 32'h573AFC6F;	14'h0477: data <= 32'h5708B659;	14'h0478: data <= 32'h56D6573E;	14'h0479: data <= 32'h56A3DF2B;	14'h047A: data <= 32'h56714E31;	14'h047B: data <= 32'h563EA45D;	14'h047C: data <= 32'h560BE1BF;	14'h047D: data <= 32'h55D90663;	14'h047E: data <= 32'h55A6125A;	14'h047F: data <= 32'h557305B2;	14'h0480: data <= 32'h553FE07A;	14'h0481: data <= 32'h550CA2BF;	14'h0482: data <= 32'h54D94C92;	14'h0483: data <= 32'h54A5DE00;	14'h0484: data <= 32'h54725719;	14'h0485: data <= 32'h543EB7EB;	14'h0486: data <= 32'h540B0085;	14'h0487: data <= 32'h53D730F6;	14'h0488: data <= 32'h53A3494D;	14'h0489: data <= 32'h536F4999;	14'h048A: data <= 32'h533B31E9;	14'h048B: data <= 32'h5307024B;	14'h048C: data <= 32'h52D2BAD0;	14'h048D: data <= 32'h529E5B85;	14'h048E: data <= 32'h5269E47A;	14'h048F: data <= 32'h523555BD;	14'h0490: data <= 32'h5200AF5F;	14'h0491: data <= 32'h51CBF16E;	14'h0492: data <= 32'h51971BFA;	14'h0493: data <= 32'h51622F11;	14'h0494: data <= 32'h512D2AC2;	14'h0495: data <= 32'h50F80F1E;	14'h0496: data <= 32'h50C2DC33;	14'h0497: data <= 32'h508D9210;	14'h0498: data <= 32'h505830C5;	14'h0499: data <= 32'h5022B862;	14'h049A: data <= 32'h4FED28F5;	14'h049B: data <= 32'h4FB7828E;	14'h049C: data <= 32'h4F81C53C;	14'h049D: data <= 32'h4F4BF10F;	14'h049E: data <= 32'h4F160617;	14'h049F: data <= 32'h4EE00462;	14'h04A0: data <= 32'h4EA9EC01;	14'h04A1: data <= 32'h4E73BD02;	14'h04A2: data <= 32'h4E3D7776;	14'h04A3: data <= 32'h4E071B6D;	14'h04A4: data <= 32'h4DD0A8F4;	14'h04A5: data <= 32'h4D9A201D;	14'h04A6: data <= 32'h4D6380F8;	14'h04A7: data <= 32'h4D2CCB93;	14'h04A8: data <= 32'h4CF5FFFE;	14'h04A9: data <= 32'h4CBF1E4A;	14'h04AA: data <= 32'h4C882685;	14'h04AB: data <= 32'h4C5118C0;	14'h04AC: data <= 32'h4C19F50B;	14'h04AD: data <= 32'h4BE2BB76;	14'h04AE: data <= 32'h4BAB6C10;	14'h04AF: data <= 32'h4B7406E9;	14'h04B0: data <= 32'h4B3C8C11;	14'h04B1: data <= 32'h4B04FB98;	14'h04B2: data <= 32'h4ACD558E;	14'h04B3: data <= 32'h4A959A04;	14'h04B4: data <= 32'h4A5DC908;	14'h04B5: data <= 32'h4A25E2AC;	14'h04B6: data <= 32'h49EDE6FF;	14'h04B7: data <= 32'h49B5D611;	14'h04B8: data <= 32'h497DAFF3;	14'h04B9: data <= 32'h494574B4;	14'h04BA: data <= 32'h490D2465;	14'h04BB: data <= 32'h48D4BF16;	14'h04BC: data <= 32'h489C44D7;	14'h04BD: data <= 32'h4863B5B9;	14'h04BE: data <= 32'h482B11CB;	14'h04BF: data <= 32'h47F2591E;	14'h04C0: data <= 32'h47B98BC2;	14'h04C1: data <= 32'h4780A9C8;	14'h04C2: data <= 32'h4747B33F;	14'h04C3: data <= 32'h470EA839;	14'h04C4: data <= 32'h46D588C6;	14'h04C5: data <= 32'h469C54F6;	14'h04C6: data <= 32'h46630CD9;	14'h04C7: data <= 32'h4629B080;	14'h04C8: data <= 32'h45F03FFC;	14'h04C9: data <= 32'h45B6BB5D;	14'h04CA: data <= 32'h457D22B3;	14'h04CB: data <= 32'h4543760F;	14'h04CC: data <= 32'h4509B583;	14'h04CD: data <= 32'h44CFE11D;	14'h04CE: data <= 32'h4495F8EF;	14'h04CF: data <= 32'h445BFD0A;	14'h04D0: data <= 32'h4421ED7E;	14'h04D1: data <= 32'h43E7CA5C;	14'h04D2: data <= 32'h43AD93B5;	14'h04D3: data <= 32'h43734999;	14'h04D4: data <= 32'h4338EC19;	14'h04D5: data <= 32'h42FE7B46;	14'h04D6: data <= 32'h42C3F731;	14'h04D7: data <= 32'h42895FEA;	14'h04D8: data <= 32'h424EB583;	14'h04D9: data <= 32'h4213F80C;	14'h04DA: data <= 32'h41D92796;	14'h04DB: data <= 32'h419E4432;	14'h04DC: data <= 32'h41634DF1;	14'h04DD: data <= 32'h412844E3;	14'h04DE: data <= 32'h40ED291B;	14'h04DF: data <= 32'h40B1FAA9;	14'h04E0: data <= 32'h4076B99D;	14'h04E1: data <= 32'h403B660A;	14'h04E2: data <= 32'h3FFFFFFF;	14'h04E3: data <= 32'h3FC4878E;	14'h04E4: data <= 32'h3F88FCC9;	14'h04E5: data <= 32'h3F4D5FC0;	14'h04E6: data <= 32'h3F11B084;	14'h04E7: data <= 32'h3ED5EF27;	14'h04E8: data <= 32'h3E9A1BB9;	14'h04E9: data <= 32'h3E5E364C;	14'h04EA: data <= 32'h3E223EF2;	14'h04EB: data <= 32'h3DE635BB;	14'h04EC: data <= 32'h3DAA1AB9;	14'h04ED: data <= 32'h3D6DEDFC;	14'h04EE: data <= 32'h3D31AF97;	14'h04EF: data <= 32'h3CF55F9A;	14'h04F0: data <= 32'h3CB8FE17;	14'h04F1: data <= 32'h3C7C8B1F;	14'h04F2: data <= 32'h3C4006C4;	14'h04F3: data <= 32'h3C037117;	14'h04F4: data <= 32'h3BC6CA2A;	14'h04F5: data <= 32'h3B8A120D;	14'h04F6: data <= 32'h3B4D48D3;	14'h04F7: data <= 32'h3B106E8C;	14'h04F8: data <= 32'h3AD3834B;	14'h04F9: data <= 32'h3A968720;	14'h04FA: data <= 32'h3A597A1E;	14'h04FB: data <= 32'h3A1C5C56;	14'h04FC: data <= 32'h39DF2DD9;	14'h04FD: data <= 32'h39A1EEB9;	14'h04FE: data <= 32'h39649F08;	14'h04FF: data <= 32'h39273ED7;	14'h0500: data <= 32'h38E9CE38;	14'h0501: data <= 32'h38AC4D3C;	14'h0502: data <= 32'h386EBBF6;	14'h0503: data <= 32'h38311A77;	14'h0504: data <= 32'h37F368D0;	14'h0505: data <= 32'h37B5A714;	14'h0506: data <= 32'h3777D554;	14'h0507: data <= 32'h3739F3A2;	14'h0508: data <= 32'h36FC0210;	14'h0509: data <= 32'h36BE00AF;	14'h050A: data <= 32'h367FEF91;	14'h050B: data <= 32'h3641CEC9;	14'h050C: data <= 32'h36039E68;	14'h050D: data <= 32'h35C55E80;	14'h050E: data <= 32'h35870F22;	14'h050F: data <= 32'h3548B061;	14'h0510: data <= 32'h350A424F;	14'h0511: data <= 32'h34CBC4FE;	14'h0512: data <= 32'h348D387F;	14'h0513: data <= 32'h344E9CE5;	14'h0514: data <= 32'h340FF241;	14'h0515: data <= 32'h33D138A6;	14'h0516: data <= 32'h33927025;	14'h0517: data <= 32'h335398D2;	14'h0518: data <= 32'h3314B2BC;	14'h0519: data <= 32'h32D5BDF8;	14'h051A: data <= 32'h3296BA97;	14'h051B: data <= 32'h3257A8AA;	14'h051C: data <= 32'h32188845;	14'h051D: data <= 32'h31D95979;	14'h051E: data <= 32'h319A1C58;	14'h051F: data <= 32'h315AD0F5;	14'h0520: data <= 32'h311B7762;	14'h0521: data <= 32'h30DC0FB1;	14'h0522: data <= 32'h309C99F5;	14'h0523: data <= 32'h305D163E;	14'h0524: data <= 32'h301D84A1;	14'h0525: data <= 32'h2FDDE52E;	14'h0526: data <= 32'h2F9E37F9;	14'h0527: data <= 32'h2F5E7D14;	14'h0528: data <= 32'h2F1EB490;	14'h0529: data <= 32'h2EDEDE81;	14'h052A: data <= 32'h2E9EFAF9;	14'h052B: data <= 32'h2E5F0A09;	14'h052C: data <= 32'h2E1F0BC5;	14'h052D: data <= 32'h2DDF003F;	14'h052E: data <= 32'h2D9EE789;	14'h052F: data <= 32'h2D5EC1B5;	14'h0530: data <= 32'h2D1E8ED7;	14'h0531: data <= 32'h2CDE4F00;	14'h0532: data <= 32'h2C9E0243;	14'h0533: data <= 32'h2C5DA8B3;	14'h0534: data <= 32'h2C1D4261;	14'h0535: data <= 32'h2BDCCF61;	14'h0536: data <= 32'h2B9C4FC5;	14'h0537: data <= 32'h2B5BC3A0;	14'h0538: data <= 32'h2B1B2B04;	14'h0539: data <= 32'h2ADA8603;	14'h053A: data <= 32'h2A99D4B1;	14'h053B: data <= 32'h2A59171F;	14'h053C: data <= 32'h2A184D61;	14'h053D: data <= 32'h29D7778A;	14'h053E: data <= 32'h299695AA;	14'h053F: data <= 32'h2955A7D7;	14'h0540: data <= 32'h2914AE21;	14'h0541: data <= 32'h28D3A89C;	14'h0542: data <= 32'h2892975B;	14'h0543: data <= 32'h28517A6F;	14'h0544: data <= 32'h281051ED;	14'h0545: data <= 32'h27CF1DE6;	14'h0546: data <= 32'h278DDE6E;	14'h0547: data <= 32'h274C9396;	14'h0548: data <= 32'h270B3D72;	14'h0549: data <= 32'h26C9DC16;	14'h054A: data <= 32'h26886F92;	14'h054B: data <= 32'h2646F7FB;	14'h054C: data <= 32'h26057562;	14'h054D: data <= 32'h25C3E7DC;	14'h054E: data <= 32'h25824F7A;	14'h054F: data <= 32'h2540AC50;	14'h0550: data <= 32'h24FEFE71;	14'h0551: data <= 32'h24BD45EF;	14'h0552: data <= 32'h247B82DD;	14'h0553: data <= 32'h2439B54E;	14'h0554: data <= 32'h23F7DD55;	14'h0555: data <= 32'h23B5FB05;	14'h0556: data <= 32'h23740E72;	14'h0557: data <= 32'h233217AD;	14'h0558: data <= 32'h22F016C9;	14'h0559: data <= 32'h22AE0BDB;	14'h055A: data <= 32'h226BF6F5;	14'h055B: data <= 32'h2229D829;	14'h055C: data <= 32'h21E7AF8B;	14'h055D: data <= 32'h21A57D2E;	14'h055E: data <= 32'h21634125;	14'h055F: data <= 32'h2120FB82;	14'h0560: data <= 32'h20DEAC5A;	14'h0561: data <= 32'h209C53BF;	14'h0562: data <= 32'h2059F1C3;	14'h0563: data <= 32'h2017867B;	14'h0564: data <= 32'h1FD511F9;	14'h0565: data <= 32'h1F929451;	14'h0566: data <= 32'h1F500D95;	14'h0567: data <= 32'h1F0D7DD8;	14'h0568: data <= 32'h1ECAE52F;	14'h0569: data <= 32'h1E8843AB;	14'h056A: data <= 32'h1E459960;	14'h056B: data <= 32'h1E02E662;	14'h056C: data <= 32'h1DC02AC2;	14'h056D: data <= 32'h1D7D6696;	14'h056E: data <= 32'h1D3A99EF;	14'h056F: data <= 32'h1CF7C4E1;	14'h0570: data <= 32'h1CB4E77F;	14'h0571: data <= 32'h1C7201DD;	14'h0572: data <= 32'h1C2F140D;	14'h0573: data <= 32'h1BEC1E23;	14'h0574: data <= 32'h1BA92032;	14'h0575: data <= 32'h1B661A4E;	14'h0576: data <= 32'h1B230C89;	14'h0577: data <= 32'h1ADFF6F7;	14'h0578: data <= 32'h1A9CD9AC;	14'h0579: data <= 32'h1A59B4B9;	14'h057A: data <= 32'h1A168834;	14'h057B: data <= 32'h19D3542F;	14'h057C: data <= 32'h199018BD;	14'h057D: data <= 32'h194CD5F2;	14'h057E: data <= 32'h19098BE1;	14'h057F: data <= 32'h18C63A9D;	14'h0580: data <= 32'h1882E23A;	14'h0581: data <= 32'h183F82CC;	14'h0582: data <= 32'h17FC1C64;	14'h0583: data <= 32'h17B8AF18;	14'h0584: data <= 32'h17753AFA;	14'h0585: data <= 32'h1731C01E;	14'h0586: data <= 32'h16EE3E96;	14'h0587: data <= 32'h16AAB677;	14'h0588: data <= 32'h166727D4;	14'h0589: data <= 32'h162392C1;	14'h058A: data <= 32'h15DFF750;	14'h058B: data <= 32'h159C5595;	14'h058C: data <= 32'h1558ADA4;	14'h058D: data <= 32'h1514FF90;	14'h058E: data <= 32'h14D14B6C;	14'h058F: data <= 32'h148D914D;	14'h0590: data <= 32'h1449D144;	14'h0591: data <= 32'h14060B67;	14'h0592: data <= 32'h13C23FC8;	14'h0593: data <= 32'h137E6E7B;	14'h0594: data <= 32'h133A9793;	14'h0595: data <= 32'h12F6BB25;	14'h0596: data <= 32'h12B2D942;	14'h0597: data <= 32'h126EF200;	14'h0598: data <= 32'h122B0571;	14'h0599: data <= 32'h11E713A9;	14'h059A: data <= 32'h11A31CBB;	14'h059B: data <= 32'h115F20BC;	14'h059C: data <= 32'h111B1FBE;	14'h059D: data <= 32'h10D719D5;	14'h059E: data <= 32'h10930F15;	14'h059F: data <= 32'h104EFF91;	14'h05A0: data <= 32'h100AEB5D;	14'h05A1: data <= 32'h0FC6D28C;	14'h05A2: data <= 32'h0F82B532;	14'h05A3: data <= 32'h0F3E9363;	14'h05A4: data <= 32'h0EFA6D32;	14'h05A5: data <= 32'h0EB642B3;	14'h05A6: data <= 32'h0E7213F8;	14'h05A7: data <= 32'h0E2DE117;	14'h05A8: data <= 32'h0DE9AA23;	14'h05A9: data <= 32'h0DA56F2E;	14'h05AA: data <= 32'h0D61304D;	14'h05AB: data <= 32'h0D1CED93;	14'h05AC: data <= 32'h0CD8A715;	14'h05AD: data <= 32'h0C945CE5;	14'h05AE: data <= 32'h0C500F17;	14'h05AF: data <= 32'h0C0BBDBF;	14'h05B0: data <= 32'h0BC768F1;	14'h05B1: data <= 32'h0B8310C0;	14'h05B2: data <= 32'h0B3EB53F;	14'h05B3: data <= 32'h0AFA5684;	14'h05B4: data <= 32'h0AB5F4A0;	14'h05B5: data <= 32'h0A718FA8;	14'h05B6: data <= 32'h0A2D27AF;	14'h05B7: data <= 32'h09E8BCC9;	14'h05B8: data <= 32'h09A44F0B;	14'h05B9: data <= 32'h095FDE86;	14'h05BA: data <= 32'h091B6B50;	14'h05BB: data <= 32'h08D6F57B;	14'h05BC: data <= 32'h08927D1C;	14'h05BD: data <= 32'h084E0246;	14'h05BE: data <= 32'h0809850D;	14'h05BF: data <= 32'h07C50585;	14'h05C0: data <= 32'h078083C0;	14'h05C1: data <= 32'h073BFFD4;	14'h05C2: data <= 32'h06F779D3;	14'h05C3: data <= 32'h06B2F1D2;	14'h05C4: data <= 32'h066E67E3;	14'h05C5: data <= 32'h0629DC1B;	14'h05C6: data <= 32'h05E54E8E;	14'h05C7: data <= 32'h05A0BF4F;	14'h05C8: data <= 32'h055C2E71;	14'h05C9: data <= 32'h05179C09;	14'h05CA: data <= 32'h04D3082A;	14'h05CB: data <= 32'h048E72E9;	14'h05CC: data <= 32'h0449DC58;	14'h05CD: data <= 32'h0405448B;	14'h05CE: data <= 32'h03C0AB96;	14'h05CF: data <= 32'h037C118E;	14'h05D0: data <= 32'h03377685;	14'h05D1: data <= 32'h02F2DA8F;	14'h05D2: data <= 32'h02AE3DC0;	14'h05D3: data <= 32'h0269A02C;	14'h05D4: data <= 32'h022501E6;	14'h05D5: data <= 32'h01E06302;	14'h05D6: data <= 32'h019BC395;	14'h05D7: data <= 32'h015723B1;	14'h05D8: data <= 32'h0112836A;	14'h05D9: data <= 32'h00CDE2D4;	14'h05DA: data <= 32'h00894204;	14'h05DB: data <= 32'h0044A10B;	14'h05DC: data <= 32'h00000000;	14'h05DD: data <= 32'hFFBB5EF5;	14'h05DE: data <= 32'hFF76BDFC;	14'h05DF: data <= 32'hFF321D2C;	14'h05E0: data <= 32'hFEED7C96;	14'h05E1: data <= 32'hFEA8DC4F;	14'h05E2: data <= 32'hFE643C6B;	14'h05E3: data <= 32'hFE1F9CFE;	14'h05E4: data <= 32'hFDDAFE1A;	14'h05E5: data <= 32'hFD965FD4;	14'h05E6: data <= 32'hFD51C240;	14'h05E7: data <= 32'hFD0D2571;	14'h05E8: data <= 32'hFCC8897B;	14'h05E9: data <= 32'hFC83EE72;	14'h05EA: data <= 32'hFC3F546A;	14'h05EB: data <= 32'hFBFABB75;	14'h05EC: data <= 32'hFBB623A8;	14'h05ED: data <= 32'hFB718D17;	14'h05EE: data <= 32'hFB2CF7D6;	14'h05EF: data <= 32'hFAE863F7;	14'h05F0: data <= 32'hFAA3D18F;	14'h05F1: data <= 32'hFA5F40B1;	14'h05F2: data <= 32'hFA1AB172;	14'h05F3: data <= 32'hF9D623E5;	14'h05F4: data <= 32'hF991981D;	14'h05F5: data <= 32'hF94D0E2E;	14'h05F6: data <= 32'hF908862D;	14'h05F7: data <= 32'hF8C4002C;	14'h05F8: data <= 32'hF87F7C40;	14'h05F9: data <= 32'hF83AFA7B;	14'h05FA: data <= 32'hF7F67AF3;	14'h05FB: data <= 32'hF7B1FDBA;	14'h05FC: data <= 32'hF76D82E4;	14'h05FD: data <= 32'hF7290A85;	14'h05FE: data <= 32'hF6E494B0;	14'h05FF: data <= 32'hF6A0217A;	14'h0600: data <= 32'hF65BB0F5;	14'h0601: data <= 32'hF6174337;	14'h0602: data <= 32'hF5D2D851;	14'h0603: data <= 32'hF58E7058;	14'h0604: data <= 32'hF54A0B60;	14'h0605: data <= 32'hF505A97C;	14'h0606: data <= 32'hF4C14AC1;	14'h0607: data <= 32'hF47CEF40;	14'h0608: data <= 32'hF438970F;	14'h0609: data <= 32'hF3F44241;	14'h060A: data <= 32'hF3AFF0E9;	14'h060B: data <= 32'hF36BA31B;	14'h060C: data <= 32'hF32758EB;	14'h060D: data <= 32'hF2E3126D;	14'h060E: data <= 32'hF29ECFB3;	14'h060F: data <= 32'hF25A90D2;	14'h0610: data <= 32'hF21655DD;	14'h0611: data <= 32'hF1D21EE9;	14'h0612: data <= 32'hF18DEC08;	14'h0613: data <= 32'hF149BD4D;	14'h0614: data <= 32'hF10592CE;	14'h0615: data <= 32'hF0C16C9D;	14'h0616: data <= 32'hF07D4ACE;	14'h0617: data <= 32'hF0392D74;	14'h0618: data <= 32'hEFF514A3;	14'h0619: data <= 32'hEFB1006F;	14'h061A: data <= 32'hEF6CF0EB;	14'h061B: data <= 32'hEF28E62B;	14'h061C: data <= 32'hEEE4E042;	14'h061D: data <= 32'hEEA0DF44;	14'h061E: data <= 32'hEE5CE345;	14'h061F: data <= 32'hEE18EC57;	14'h0620: data <= 32'hEDD4FA8F;	14'h0621: data <= 32'hED910E00;	14'h0622: data <= 32'hED4D26BE;	14'h0623: data <= 32'hED0944DB;	14'h0624: data <= 32'hECC5686D;	14'h0625: data <= 32'hEC819185;	14'h0626: data <= 32'hEC3DC038;	14'h0627: data <= 32'hEBF9F499;	14'h0628: data <= 32'hEBB62EBC;	14'h0629: data <= 32'hEB726EB3;	14'h062A: data <= 32'hEB2EB494;	14'h062B: data <= 32'hEAEB0070;	14'h062C: data <= 32'hEAA7525C;	14'h062D: data <= 32'hEA63AA6B;	14'h062E: data <= 32'hEA2008B0;	14'h062F: data <= 32'hE9DC6D3F;	14'h0630: data <= 32'hE998D82C;	14'h0631: data <= 32'hE9554989;	14'h0632: data <= 32'hE911C16A;	14'h0633: data <= 32'hE8CE3FE2;	14'h0634: data <= 32'hE88AC506;	14'h0635: data <= 32'hE84750E8;	14'h0636: data <= 32'hE803E39C;	14'h0637: data <= 32'hE7C07D34;	14'h0638: data <= 32'hE77D1DC6;	14'h0639: data <= 32'hE739C563;	14'h063A: data <= 32'hE6F6741F;	14'h063B: data <= 32'hE6B32A0E;	14'h063C: data <= 32'hE66FE743;	14'h063D: data <= 32'hE62CABD1;	14'h063E: data <= 32'hE5E977CC;	14'h063F: data <= 32'hE5A64B47;	14'h0640: data <= 32'hE5632654;	14'h0641: data <= 32'hE5200909;	14'h0642: data <= 32'hE4DCF377;	14'h0643: data <= 32'hE499E5B2;	14'h0644: data <= 32'hE456DFCE;	14'h0645: data <= 32'hE413E1DD;	14'h0646: data <= 32'hE3D0EBF3;	14'h0647: data <= 32'hE38DFE23;	14'h0648: data <= 32'hE34B1881;	14'h0649: data <= 32'hE3083B1F;	14'h064A: data <= 32'hE2C56611;	14'h064B: data <= 32'hE282996A;	14'h064C: data <= 32'hE23FD53E;	14'h064D: data <= 32'hE1FD199E;	14'h064E: data <= 32'hE1BA66A0;	14'h064F: data <= 32'hE177BC55;	14'h0650: data <= 32'hE1351AD1;	14'h0651: data <= 32'hE0F28228;	14'h0652: data <= 32'hE0AFF26B;	14'h0653: data <= 32'hE06D6BAF;	14'h0654: data <= 32'hE02AEE07;	14'h0655: data <= 32'hDFE87985;	14'h0656: data <= 32'hDFA60E3D;	14'h0657: data <= 32'hDF63AC41;	14'h0658: data <= 32'hDF2153A6;	14'h0659: data <= 32'hDEDF047E;	14'h065A: data <= 32'hDE9CBEDB;	14'h065B: data <= 32'hDE5A82D2;	14'h065C: data <= 32'hDE185075;	14'h065D: data <= 32'hDDD627D7;	14'h065E: data <= 32'hDD94090B;	14'h065F: data <= 32'hDD51F425;	14'h0660: data <= 32'hDD0FE937;	14'h0661: data <= 32'hDCCDE853;	14'h0662: data <= 32'hDC8BF18E;	14'h0663: data <= 32'hDC4A04FB;	14'h0664: data <= 32'hDC0822AB;	14'h0665: data <= 32'hDBC64AB2;	14'h0666: data <= 32'hDB847D23;	14'h0667: data <= 32'hDB42BA11;	14'h0668: data <= 32'hDB01018F;	14'h0669: data <= 32'hDABF53B0;	14'h066A: data <= 32'hDA7DB086;	14'h066B: data <= 32'hDA3C1824;	14'h066C: data <= 32'hD9FA8A9E;	14'h066D: data <= 32'hD9B90805;	14'h066E: data <= 32'hD977906E;	14'h066F: data <= 32'hD93623EA;	14'h0670: data <= 32'hD8F4C28E;	14'h0671: data <= 32'hD8B36C6A;	14'h0672: data <= 32'hD8722192;	14'h0673: data <= 32'hD830E21A;	14'h0674: data <= 32'hD7EFAE13;	14'h0675: data <= 32'hD7AE8591;	14'h0676: data <= 32'hD76D68A5;	14'h0677: data <= 32'hD72C5764;	14'h0678: data <= 32'hD6EB51DF;	14'h0679: data <= 32'hD6AA5829;	14'h067A: data <= 32'hD6696A56;	14'h067B: data <= 32'hD6288876;	14'h067C: data <= 32'hD5E7B29F;	14'h067D: data <= 32'hD5A6E8E1;	14'h067E: data <= 32'hD5662B4F;	14'h067F: data <= 32'hD52579FD;	14'h0680: data <= 32'hD4E4D4FC;	14'h0681: data <= 32'hD4A43C60;	14'h0682: data <= 32'hD463B03B;	14'h0683: data <= 32'hD423309F;	14'h0684: data <= 32'hD3E2BD9F;	14'h0685: data <= 32'hD3A2574D;	14'h0686: data <= 32'hD361FDBD;	14'h0687: data <= 32'hD321B100;	14'h0688: data <= 32'hD2E17129;	14'h0689: data <= 32'hD2A13E4B;	14'h068A: data <= 32'hD2611877;	14'h068B: data <= 32'hD220FFC1;	14'h068C: data <= 32'hD1E0F43B;	14'h068D: data <= 32'hD1A0F5F7;	14'h068E: data <= 32'hD1610507;	14'h068F: data <= 32'hD121217F;	14'h0690: data <= 32'hD0E14B70;	14'h0691: data <= 32'hD0A182EC;	14'h0692: data <= 32'hD061C807;	14'h0693: data <= 32'hD0221AD2;	14'h0694: data <= 32'hCFE27B5F;	14'h0695: data <= 32'hCFA2E9C2;	14'h0696: data <= 32'hCF63660B;	14'h0697: data <= 32'hCF23F04F;	14'h0698: data <= 32'hCEE4889E;	14'h0699: data <= 32'hCEA52F0B;	14'h069A: data <= 32'hCE65E3A8;	14'h069B: data <= 32'hCE26A687;	14'h069C: data <= 32'hCDE777BB;	14'h069D: data <= 32'hCDA85756;	14'h069E: data <= 32'hCD694569;	14'h069F: data <= 32'hCD2A4208;	14'h06A0: data <= 32'hCCEB4D44;	14'h06A1: data <= 32'hCCAC672E;	14'h06A2: data <= 32'hCC6D8FDB;	14'h06A3: data <= 32'hCC2EC75A;	14'h06A4: data <= 32'hCBF00DBF;	14'h06A5: data <= 32'hCBB1631B;	14'h06A6: data <= 32'hCB72C781;	14'h06A7: data <= 32'hCB343B02;	14'h06A8: data <= 32'hCAF5BDB1;	14'h06A9: data <= 32'hCAB74F9F;	14'h06AA: data <= 32'hCA78F0DE;	14'h06AB: data <= 32'hCA3AA180;	14'h06AC: data <= 32'hC9FC6198;	14'h06AD: data <= 32'hC9BE3137;	14'h06AE: data <= 32'hC980106F;	14'h06AF: data <= 32'hC941FF51;	14'h06B0: data <= 32'hC903FDF0;	14'h06B1: data <= 32'hC8C60C5E;	14'h06B2: data <= 32'hC8882AAC;	14'h06B3: data <= 32'hC84A58EC;	14'h06B4: data <= 32'hC80C9730;	14'h06B5: data <= 32'hC7CEE589;	14'h06B6: data <= 32'hC791440A;	14'h06B7: data <= 32'hC753B2C4;	14'h06B8: data <= 32'hC71631C8;	14'h06B9: data <= 32'hC6D8C129;	14'h06BA: data <= 32'hC69B60F8;	14'h06BB: data <= 32'hC65E1147;	14'h06BC: data <= 32'hC620D227;	14'h06BD: data <= 32'hC5E3A3AA;	14'h06BE: data <= 32'hC5A685E2;	14'h06BF: data <= 32'hC56978E0;	14'h06C0: data <= 32'hC52C7CB5;	14'h06C1: data <= 32'hC4EF9174;	14'h06C2: data <= 32'hC4B2B72D;	14'h06C3: data <= 32'hC475EDF3;	14'h06C4: data <= 32'hC43935D6;	14'h06C5: data <= 32'hC3FC8EE9;	14'h06C6: data <= 32'hC3BFF93C;	14'h06C7: data <= 32'hC38374E1;	14'h06C8: data <= 32'hC34701E9;	14'h06C9: data <= 32'hC30AA066;	14'h06CA: data <= 32'hC2CE5069;	14'h06CB: data <= 32'hC2921204;	14'h06CC: data <= 32'hC255E547;	14'h06CD: data <= 32'hC219CA45;	14'h06CE: data <= 32'hC1DDC10E;	14'h06CF: data <= 32'hC1A1C9B4;	14'h06D0: data <= 32'hC165E447;	14'h06D1: data <= 32'hC12A10D9;	14'h06D2: data <= 32'hC0EE4F7C;	14'h06D3: data <= 32'hC0B2A040;	14'h06D4: data <= 32'hC0770337;	14'h06D5: data <= 32'hC03B7872;	14'h06D6: data <= 32'hC0000001;	14'h06D7: data <= 32'hBFC499F6;	14'h06D8: data <= 32'hBF894663;	14'h06D9: data <= 32'hBF4E0557;	14'h06DA: data <= 32'hBF12D6E5;	14'h06DB: data <= 32'hBED7BB1D;	14'h06DC: data <= 32'hBE9CB20F;	14'h06DD: data <= 32'hBE61BBCE;	14'h06DE: data <= 32'hBE26D86A;	14'h06DF: data <= 32'hBDEC07F4;	14'h06E0: data <= 32'hBDB14A7D;	14'h06E1: data <= 32'hBD76A016;	14'h06E2: data <= 32'hBD3C08CF;	14'h06E3: data <= 32'hBD0184BA;	14'h06E4: data <= 32'hBCC713E7;	14'h06E5: data <= 32'hBC8CB667;	14'h06E6: data <= 32'hBC526C4B;	14'h06E7: data <= 32'hBC1835A4;	14'h06E8: data <= 32'hBBDE1282;	14'h06E9: data <= 32'hBBA402F6;	14'h06EA: data <= 32'hBB6A0711;	14'h06EB: data <= 32'hBB301EE3;	14'h06EC: data <= 32'hBAF64A7D;	14'h06ED: data <= 32'hBABC89F1;	14'h06EE: data <= 32'hBA82DD4D;	14'h06EF: data <= 32'hBA4944A3;	14'h06F0: data <= 32'hBA0FC004;	14'h06F1: data <= 32'hB9D64F80;	14'h06F2: data <= 32'hB99CF327;	14'h06F3: data <= 32'hB963AB0A;	14'h06F4: data <= 32'hB92A773A;	14'h06F5: data <= 32'hB8F157C7;	14'h06F6: data <= 32'hB8B84CC1;	14'h06F7: data <= 32'hB87F5638;	14'h06F8: data <= 32'hB846743E;	14'h06F9: data <= 32'hB80DA6E2;	14'h06FA: data <= 32'hB7D4EE35;	14'h06FB: data <= 32'hB79C4A47;	14'h06FC: data <= 32'hB763BB29;	14'h06FD: data <= 32'hB72B40EA;	14'h06FE: data <= 32'hB6F2DB9B;	14'h06FF: data <= 32'hB6BA8B4C;	14'h0700: data <= 32'hB682500D;	14'h0701: data <= 32'hB64A29EF;	14'h0702: data <= 32'hB6121901;	14'h0703: data <= 32'hB5DA1D54;	14'h0704: data <= 32'hB5A236F8;	14'h0705: data <= 32'hB56A65FC;	14'h0706: data <= 32'hB532AA72;	14'h0707: data <= 32'hB4FB0468;	14'h0708: data <= 32'hB4C373EF;	14'h0709: data <= 32'hB48BF917;	14'h070A: data <= 32'hB45493F0;	14'h070B: data <= 32'hB41D448A;	14'h070C: data <= 32'hB3E60AF5;	14'h070D: data <= 32'hB3AEE740;	14'h070E: data <= 32'hB377D97B;	14'h070F: data <= 32'hB340E1B6;	14'h0710: data <= 32'hB30A0002;	14'h0711: data <= 32'hB2D3346D;	14'h0712: data <= 32'hB29C7F08;	14'h0713: data <= 32'hB265DFE3;	14'h0714: data <= 32'hB22F570C;	14'h0715: data <= 32'hB1F8E493;	14'h0716: data <= 32'hB1C2888A;	14'h0717: data <= 32'hB18C42FE;	14'h0718: data <= 32'hB15613FF;	14'h0719: data <= 32'hB11FFB9E;	14'h071A: data <= 32'hB0E9F9E9;	14'h071B: data <= 32'hB0B40EF1;	14'h071C: data <= 32'hB07E3AC4;	14'h071D: data <= 32'hB0487D72;	14'h071E: data <= 32'hB012D70B;	14'h071F: data <= 32'hAFDD479E;	14'h0720: data <= 32'hAFA7CF3B;	14'h0721: data <= 32'hAF726DF0;	14'h0722: data <= 32'hAF3D23CD;	14'h0723: data <= 32'hAF07F0E2;	14'h0724: data <= 32'hAED2D53E;	14'h0725: data <= 32'hAE9DD0EF;	14'h0726: data <= 32'hAE68E406;	14'h0727: data <= 32'hAE340E92;	14'h0728: data <= 32'hADFF50A1;	14'h0729: data <= 32'hADCAAA43;	14'h072A: data <= 32'hAD961B86;	14'h072B: data <= 32'hAD61A47B;	14'h072C: data <= 32'hAD2D4530;	14'h072D: data <= 32'hACF8FDB5;	14'h072E: data <= 32'hACC4CE17;	14'h072F: data <= 32'hAC90B667;	14'h0730: data <= 32'hAC5CB6B3;	14'h0731: data <= 32'hAC28CF0A;	14'h0732: data <= 32'hABF4FF7B;	14'h0733: data <= 32'hABC14815;	14'h0734: data <= 32'hAB8DA8E7;	14'h0735: data <= 32'hAB5A2200;	14'h0736: data <= 32'hAB26B36E;	14'h0737: data <= 32'hAAF35D41;	14'h0738: data <= 32'hAAC01F86;	14'h0739: data <= 32'hAA8CFA4E;	14'h073A: data <= 32'hAA59EDA6;	14'h073B: data <= 32'hAA26F99D;	14'h073C: data <= 32'hA9F41E41;	14'h073D: data <= 32'hA9C15BA3;	14'h073E: data <= 32'hA98EB1CF;	14'h073F: data <= 32'hA95C20D5;	14'h0740: data <= 32'hA929A8C2;	14'h0741: data <= 32'hA8F749A7;	14'h0742: data <= 32'hA8C50391;	14'h0743: data <= 32'hA892D68E;	14'h0744: data <= 32'hA860C2AD;	14'h0745: data <= 32'hA82EC7FC;	14'h0746: data <= 32'hA7FCE68B;	14'h0747: data <= 32'hA7CB1E66;	14'h0748: data <= 32'hA7996F9D;	14'h0749: data <= 32'hA767DA3D;	14'h074A: data <= 32'hA7365E56;	14'h074B: data <= 32'hA704FBF4;	14'h074C: data <= 32'hA6D3B327;	14'h074D: data <= 32'hA6A283FC;	14'h074E: data <= 32'hA6716E82;	14'h074F: data <= 32'hA64072C7;	14'h0750: data <= 32'hA60F90D9;	14'h0751: data <= 32'hA5DEC8C5;	14'h0752: data <= 32'hA5AE1A9B;	14'h0753: data <= 32'hA57D8667;	14'h0754: data <= 32'hA54D0C39;	14'h0755: data <= 32'hA51CAC1D;	14'h0756: data <= 32'hA4EC6621;	14'h0757: data <= 32'hA4BC3A55;	14'h0758: data <= 32'hA48C28C5;	14'h0759: data <= 32'hA45C317F;	14'h075A: data <= 32'hA42C5491;	14'h075B: data <= 32'hA3FC9209;	14'h075C: data <= 32'hA3CCE9F5;	14'h075D: data <= 32'hA39D5C62;	14'h075E: data <= 32'hA36DE95D;	14'h075F: data <= 32'hA33E90F6;	14'h0760: data <= 32'hA30F5338;	14'h0761: data <= 32'hA2E03032;	14'h0762: data <= 32'hA2B127F2;	14'h0763: data <= 32'hA2823A84;	14'h0764: data <= 32'hA25367F7;	14'h0765: data <= 32'hA224B057;	14'h0766: data <= 32'hA1F613B3;	14'h0767: data <= 32'hA1C79217;	14'h0768: data <= 32'hA1992B92;	14'h0769: data <= 32'hA16AE02F;	14'h076A: data <= 32'hA13CAFFD;	14'h076B: data <= 32'hA10E9B09;	14'h076C: data <= 32'hA0E0A160;	14'h076D: data <= 32'hA0B2C310;	14'h076E: data <= 32'hA0850025;	14'h076F: data <= 32'hA05758AD;	14'h0770: data <= 32'hA029CCB4;	14'h0771: data <= 32'h9FFC5C49;	14'h0772: data <= 32'h9FCF0778;	14'h0773: data <= 32'h9FA1CE4D;	14'h0774: data <= 32'h9F74B0D7;	14'h0775: data <= 32'h9F47AF21;	14'h0776: data <= 32'h9F1AC93A;	14'h0777: data <= 32'h9EEDFF2D;	14'h0778: data <= 32'h9EC15108;	14'h0779: data <= 32'h9E94BED7;	14'h077A: data <= 32'h9E6848A8;	14'h077B: data <= 32'h9E3BEE87;	14'h077C: data <= 32'h9E0FB081;	14'h077D: data <= 32'h9DE38EA3;	14'h077E: data <= 32'h9DB788F9;	14'h077F: data <= 32'h9D8B9F8F;	14'h0780: data <= 32'h9D5FD274;	14'h0781: data <= 32'h9D3421B2;	14'h0782: data <= 32'h9D088D58;	14'h0783: data <= 32'h9CDD1570;	14'h0784: data <= 32'h9CB1BA08;	14'h0785: data <= 32'h9C867B2D;	14'h0786: data <= 32'h9C5B58EA;	14'h0787: data <= 32'h9C30534C;	14'h0788: data <= 32'h9C056A60;	14'h0789: data <= 32'h9BDA9E31;	14'h078A: data <= 32'h9BAFEECD;	14'h078B: data <= 32'h9B855C3E;	14'h078C: data <= 32'h9B5AE693;	14'h078D: data <= 32'h9B308DD6;	14'h078E: data <= 32'h9B065214;	14'h078F: data <= 32'h9ADC3359;	14'h0790: data <= 32'h9AB231B1;	14'h0791: data <= 32'h9A884D29;	14'h0792: data <= 32'h9A5E85CC;	14'h0793: data <= 32'h9A34DBA6;	14'h0794: data <= 32'h9A0B4EC3;	14'h0795: data <= 32'h99E1DF30;	14'h0796: data <= 32'h99B88CF8;	14'h0797: data <= 32'h998F5827;	14'h0798: data <= 32'h996640C9;	14'h0799: data <= 32'h993D46E9;	14'h079A: data <= 32'h99146A94;	14'h079B: data <= 32'h98EBABD5;	14'h079C: data <= 32'h98C30AB8;	14'h079D: data <= 32'h989A8749;	14'h079E: data <= 32'h98722193;	14'h079F: data <= 32'h9849D9A2;	14'h07A0: data <= 32'h9821AF81;	14'h07A1: data <= 32'h97F9A33C;	14'h07A2: data <= 32'h97D1B4DF;	14'h07A3: data <= 32'h97A9E475;	14'h07A4: data <= 32'h97823209;	14'h07A5: data <= 32'h975A9DA7;	14'h07A6: data <= 32'h9733275B;	14'h07A7: data <= 32'h970BCF2E;	14'h07A8: data <= 32'h96E4952E;	14'h07A9: data <= 32'h96BD7965;	14'h07AA: data <= 32'h96967BDE;	14'h07AB: data <= 32'h966F9CA5;	14'h07AC: data <= 32'h9648DBC5;	14'h07AD: data <= 32'h96223948;	14'h07AE: data <= 32'h95FBB53B;	14'h07AF: data <= 32'h95D54FA8;	14'h07B0: data <= 32'h95AF089A;	14'h07B1: data <= 32'h9588E01C;	14'h07B2: data <= 32'h9562D639;	14'h07B3: data <= 32'h953CEAFC;	14'h07B4: data <= 32'h95171E70;	14'h07B5: data <= 32'h94F170A0;	14'h07B6: data <= 32'h94CBE197;	14'h07B7: data <= 32'h94A6715F;	14'h07B8: data <= 32'h94812003;	14'h07B9: data <= 32'h945BED8E;	14'h07BA: data <= 32'h9436DA0B;	14'h07BB: data <= 32'h9411E584;	14'h07BC: data <= 32'h93ED1004;	14'h07BD: data <= 32'h93C85995;	14'h07BE: data <= 32'h93A3C243;	14'h07BF: data <= 32'h937F4A17;	14'h07C0: data <= 32'h935AF11C;	14'h07C1: data <= 32'h9336B75D;	14'h07C2: data <= 32'h93129CE3;	14'h07C3: data <= 32'h92EEA1BA;	14'h07C4: data <= 32'h92CAC5EB;	14'h07C5: data <= 32'h92A70982;	14'h07C6: data <= 32'h92836C88;	14'h07C7: data <= 32'h925FEF07;	14'h07C8: data <= 32'h923C9109;	14'h07C9: data <= 32'h9219529A;	14'h07CA: data <= 32'h91F633C3;	14'h07CB: data <= 32'h91D3348D;	14'h07CC: data <= 32'h91B05504;	14'h07CD: data <= 32'h918D9531;	14'h07CE: data <= 32'h916AF51E;	14'h07CF: data <= 32'h914874D5;	14'h07D0: data <= 32'h91261460;	14'h07D1: data <= 32'h9103D3C9;	14'h07D2: data <= 32'h90E1B31A;	14'h07D3: data <= 32'h90BFB25C;	14'h07D4: data <= 32'h909DD199;	14'h07D5: data <= 32'h907C10DC;	14'h07D6: data <= 32'h905A702D;	14'h07D7: data <= 32'h9038EF97;	14'h07D8: data <= 32'h90178F23;	14'h07D9: data <= 32'h8FF64EDB;	14'h07DA: data <= 32'h8FD52EC7;	14'h07DB: data <= 32'h8FB42EF3;	14'h07DC: data <= 32'h8F934F66;	14'h07DD: data <= 32'h8F72902C;	14'h07DE: data <= 32'h8F51F14C;	14'h07DF: data <= 32'h8F3172D1;	14'h07E0: data <= 32'h8F1114C4;	14'h07E1: data <= 32'h8EF0D72E;	14'h07E2: data <= 32'h8ED0BA18;	14'h07E3: data <= 32'h8EB0BD8C;	14'h07E4: data <= 32'h8E90E192;	14'h07E5: data <= 32'h8E712635;	14'h07E6: data <= 32'h8E518B7C;	14'h07E7: data <= 32'h8E321172;	14'h07E8: data <= 32'h8E12B81F;	14'h07E9: data <= 32'h8DF37F8C;	14'h07EA: data <= 32'h8DD467C3;	14'h07EB: data <= 32'h8DB570CB;	14'h07EC: data <= 32'h8D969AAF;	14'h07ED: data <= 32'h8D77E577;	14'h07EE: data <= 32'h8D59512B;	14'h07EF: data <= 32'h8D3ADDD5;	14'h07F0: data <= 32'h8D1C8B7D;	14'h07F1: data <= 32'h8CFE5A2C;	14'h07F2: data <= 32'h8CE049EB;	14'h07F3: data <= 32'h8CC25AC2;	14'h07F4: data <= 32'h8CA48CBA;	14'h07F5: data <= 32'h8C86DFDB;	14'h07F6: data <= 32'h8C69542F;	14'h07F7: data <= 32'h8C4BE9BD;	14'h07F8: data <= 32'h8C2EA08E;	14'h07F9: data <= 32'h8C1178AA;	14'h07FA: data <= 32'h8BF4721B;	14'h07FB: data <= 32'h8BD78CE7;	14'h07FC: data <= 32'h8BBAC918;	14'h07FD: data <= 32'h8B9E26B5;	14'h07FE: data <= 32'h8B81A5C7;	14'h07FF: data <= 32'h8B654657;	14'h0800: data <= 32'h8B49086C;	14'h0801: data <= 32'h8B2CEC0E;	14'h0802: data <= 32'h8B10F145;	14'h0803: data <= 32'h8AF5181B;	14'h0804: data <= 32'h8AD96095;	14'h0805: data <= 32'h8ABDCABD;	14'h0806: data <= 32'h8AA2569B;	14'h0807: data <= 32'h8A870436;	14'h0808: data <= 32'h8A6BD396;	14'h0809: data <= 32'h8A50C4C3;	14'h080A: data <= 32'h8A35D7C5;	14'h080B: data <= 32'h8A1B0CA3;	14'h080C: data <= 32'h8A006366;	14'h080D: data <= 32'h89E5DC14;	14'h080E: data <= 32'h89CB76B6;	14'h080F: data <= 32'h89B13353;	14'h0810: data <= 32'h899711F3;	14'h0811: data <= 32'h897D129C;	14'h0812: data <= 32'h89633558;	14'h0813: data <= 32'h89497A2C;	14'h0814: data <= 32'h892FE121;	14'h0815: data <= 32'h89166A3E;	14'h0816: data <= 32'h88FD158A;	14'h0817: data <= 32'h88E3E30C;	14'h0818: data <= 32'h88CAD2CC;	14'h0819: data <= 32'h88B1E4D1;	14'h081A: data <= 32'h88991921;	14'h081B: data <= 32'h88806FC5;	14'h081C: data <= 32'h8867E8C4;	14'h081D: data <= 32'h884F8423;	14'h081E: data <= 32'h883741EB;	14'h081F: data <= 32'h881F2222;	14'h0820: data <= 32'h880724CF;	14'h0821: data <= 32'h87EF49FA;	14'h0822: data <= 32'h87D791A8;	14'h0823: data <= 32'h87BFFBE2;	14'h0824: data <= 32'h87A888AC;	14'h0825: data <= 32'h8791380F;	14'h0826: data <= 32'h877A0A12;	14'h0827: data <= 32'h8762FEB9;	14'h0828: data <= 32'h874C160D;	14'h0829: data <= 32'h87355014;	14'h082A: data <= 32'h871EACD5;	14'h082B: data <= 32'h87082C55;	14'h082C: data <= 32'h86F1CE9C;	14'h082D: data <= 32'h86DB93B0;	14'h082E: data <= 32'h86C57B96;	14'h082F: data <= 32'h86AF8657;	14'h0830: data <= 32'h8699B3F7;	14'h0831: data <= 32'h8684047E;	14'h0832: data <= 32'h866E77F1;	14'h0833: data <= 32'h86590E56;	14'h0834: data <= 32'h8643C7B4;	14'h0835: data <= 32'h862EA412;	14'h0836: data <= 32'h8619A374;	14'h0837: data <= 32'h8604C5E1;	14'h0838: data <= 32'h85F00B5F;	14'h0839: data <= 32'h85DB73F4;	14'h083A: data <= 32'h85C6FFA6;	14'h083B: data <= 32'h85B2AE7A;	14'h083C: data <= 32'h859E8077;	14'h083D: data <= 32'h858A75A3;	14'h083E: data <= 32'h85768E03;	14'h083F: data <= 32'h8562C99C;	14'h0840: data <= 32'h854F2875;	14'h0841: data <= 32'h853BAA94;	14'h0842: data <= 32'h85284FFD;	14'h0843: data <= 32'h851518B6;	14'h0844: data <= 32'h850204C6;	14'h0845: data <= 32'h84EF1430;	14'h0846: data <= 32'h84DC46FC;	14'h0847: data <= 32'h84C99D2E;	14'h0848: data <= 32'h84B716CB;	14'h0849: data <= 32'h84A4B3D9;	14'h084A: data <= 32'h8492745E;	14'h084B: data <= 32'h8480585D;	14'h084C: data <= 32'h846E5FDE;	14'h084D: data <= 32'h845C8AE4;	14'h084E: data <= 32'h844AD976;	14'h084F: data <= 32'h84394B97;	14'h0850: data <= 32'h8427E14D;	14'h0851: data <= 32'h84169A9E;	14'h0852: data <= 32'h8405778D;	14'h0853: data <= 32'h83F47821;	14'h0854: data <= 32'h83E39C5D;	14'h0855: data <= 32'h83D2E447;	14'h0856: data <= 32'h83C24FE4;	14'h0857: data <= 32'h83B1DF37;	14'h0858: data <= 32'h83A19247;	14'h0859: data <= 32'h83916918;	14'h085A: data <= 32'h838163AD;	14'h085B: data <= 32'h8371820D;	14'h085C: data <= 32'h8361C43C;	14'h085D: data <= 32'h83522A3D;	14'h085E: data <= 32'h8342B416;	14'h085F: data <= 32'h833361CA;	14'h0860: data <= 32'h83243360;	14'h0861: data <= 32'h831528D9;	14'h0862: data <= 32'h8306423C;	14'h0863: data <= 32'h82F77F8D;	14'h0864: data <= 32'h82E8E0CE;	14'h0865: data <= 32'h82DA6606;	14'h0866: data <= 32'h82CC0F38;	14'h0867: data <= 32'h82BDDC67;	14'h0868: data <= 32'h82AFCD99;	14'h0869: data <= 32'h82A1E2D1;	14'h086A: data <= 32'h82941C13;	14'h086B: data <= 32'h82867963;	14'h086C: data <= 32'h8278FAC6;	14'h086D: data <= 32'h826BA03E;	14'h086E: data <= 32'h825E69D0;	14'h086F: data <= 32'h82515780;	14'h0870: data <= 32'h82446951;	14'h0871: data <= 32'h82379F47;	14'h0872: data <= 32'h822AF966;	14'h0873: data <= 32'h821E77B1;	14'h0874: data <= 32'h82121A2C;	14'h0875: data <= 32'h8205E0DB;	14'h0876: data <= 32'h81F9CBC1;	14'h0877: data <= 32'h81EDDAE1;	14'h0878: data <= 32'h81E20E3F;	14'h0879: data <= 32'h81D665DF;	14'h087A: data <= 32'h81CAE1C3;	14'h087B: data <= 32'h81BF81EF;	14'h087C: data <= 32'h81B44667;	14'h087D: data <= 32'h81A92F2D;	14'h087E: data <= 32'h819E3C44;	14'h087F: data <= 32'h81936DB1;	14'h0880: data <= 32'h8188C375;	14'h0881: data <= 32'h817E3D95;	14'h0882: data <= 32'h8173DC12;	14'h0883: data <= 32'h81699EF1;	14'h0884: data <= 32'h815F8633;	14'h0885: data <= 32'h815591DC;	14'h0886: data <= 32'h814BC1EF;	14'h0887: data <= 32'h8142166F;	14'h0888: data <= 32'h81388F5E;	14'h0889: data <= 32'h812F2CBF;	14'h088A: data <= 32'h8125EE95;	14'h088B: data <= 32'h811CD4E2;	14'h088C: data <= 32'h8113DFA9;	14'h088D: data <= 32'h810B0EED;	14'h088E: data <= 32'h810262AF;	14'h088F: data <= 32'h80F9DAF4;	14'h0890: data <= 32'h80F177BD;	14'h0891: data <= 32'h80E9390C;	14'h0892: data <= 32'h80E11EE4;	14'h0893: data <= 32'h80D92947;	14'h0894: data <= 32'h80D15838;	14'h0895: data <= 32'h80C9ABB8;	14'h0896: data <= 32'h80C223CA;	14'h0897: data <= 32'h80BAC071;	14'h0898: data <= 32'h80B381AE;	14'h0899: data <= 32'h80AC6783;	14'h089A: data <= 32'h80A571F2;	14'h089B: data <= 32'h809EA0FE;	14'h089C: data <= 32'h8097F4A8;	14'h089D: data <= 32'h80916CF2;	14'h089E: data <= 32'h808B09DE;	14'h089F: data <= 32'h8084CB6F;	14'h08A0: data <= 32'h807EB1A5;	14'h08A1: data <= 32'h8078BC82;	14'h08A2: data <= 32'h8072EC09;	14'h08A3: data <= 32'h806D403B;	14'h08A4: data <= 32'h8067B919;	14'h08A5: data <= 32'h806256A5;	14'h08A6: data <= 32'h805D18E1;	14'h08A7: data <= 32'h8057FFCE;	14'h08A8: data <= 32'h80530B6D;	14'h08A9: data <= 32'h804E3BC1;	14'h08AA: data <= 32'h804990CA;	14'h08AB: data <= 32'h80450A8A;	14'h08AC: data <= 32'h8040A902;	14'h08AD: data <= 32'h803C6C33;	14'h08AE: data <= 32'h8038541F;	14'h08AF: data <= 32'h803460C7;	14'h08B0: data <= 32'h8030922B;	14'h08B1: data <= 32'h802CE84D;	14'h08B2: data <= 32'h8029632F;	14'h08B3: data <= 32'h802602D0;	14'h08B4: data <= 32'h8022C732;	14'h08B5: data <= 32'h801FB056;	14'h08B6: data <= 32'h801CBE3E;	14'h08B7: data <= 32'h8019F0E8;	14'h08B8: data <= 32'h80174857;	14'h08B9: data <= 32'h8014C48C;	14'h08BA: data <= 32'h80126586;	14'h08BB: data <= 32'h80102B47;	14'h08BC: data <= 32'h800E15CF;	14'h08BD: data <= 32'h800C251F;	14'h08BE: data <= 32'h800A5938;	14'h08BF: data <= 32'h8008B219;	14'h08C0: data <= 32'h80072FC4;	14'h08C1: data <= 32'h8005D239;	14'h08C2: data <= 32'h80049978;	14'h08C3: data <= 32'h80038581;	14'h08C4: data <= 32'h80029656;	14'h08C5: data <= 32'h8001CBF5;	14'h08C6: data <= 32'h80012660;	14'h08C7: data <= 32'h8000A597;	14'h08C8: data <= 32'h80004999;	14'h08C9: data <= 32'h80001267;	14'h08CA: data <= 32'h80000001;	14'h08CB: data <= 32'h80001267;	14'h08CC: data <= 32'h80004999;	14'h08CD: data <= 32'h8000A597;	14'h08CE: data <= 32'h80012660;	14'h08CF: data <= 32'h8001CBF5;	14'h08D0: data <= 32'h80029656;	14'h08D1: data <= 32'h80038581;	14'h08D2: data <= 32'h80049978;	14'h08D3: data <= 32'h8005D239;	14'h08D4: data <= 32'h80072FC4;	14'h08D5: data <= 32'h8008B219;	14'h08D6: data <= 32'h800A5938;	14'h08D7: data <= 32'h800C251F;	14'h08D8: data <= 32'h800E15CF;	14'h08D9: data <= 32'h80102B47;	14'h08DA: data <= 32'h80126586;	14'h08DB: data <= 32'h8014C48C;	14'h08DC: data <= 32'h80174857;	14'h08DD: data <= 32'h8019F0E8;	14'h08DE: data <= 32'h801CBE3E;	14'h08DF: data <= 32'h801FB056;	14'h08E0: data <= 32'h8022C732;	14'h08E1: data <= 32'h802602D0;	14'h08E2: data <= 32'h8029632F;	14'h08E3: data <= 32'h802CE84D;	14'h08E4: data <= 32'h8030922B;	14'h08E5: data <= 32'h803460C7;	14'h08E6: data <= 32'h8038541F;	14'h08E7: data <= 32'h803C6C33;	14'h08E8: data <= 32'h8040A902;	14'h08E9: data <= 32'h80450A8A;	14'h08EA: data <= 32'h804990CA;	14'h08EB: data <= 32'h804E3BC1;	14'h08EC: data <= 32'h80530B6D;	14'h08ED: data <= 32'h8057FFCE;	14'h08EE: data <= 32'h805D18E1;	14'h08EF: data <= 32'h806256A5;	14'h08F0: data <= 32'h8067B919;	14'h08F1: data <= 32'h806D403B;	14'h08F2: data <= 32'h8072EC09;	14'h08F3: data <= 32'h8078BC82;	14'h08F4: data <= 32'h807EB1A5;	14'h08F5: data <= 32'h8084CB6F;	14'h08F6: data <= 32'h808B09DE;	14'h08F7: data <= 32'h80916CF2;	14'h08F8: data <= 32'h8097F4A8;	14'h08F9: data <= 32'h809EA0FE;	14'h08FA: data <= 32'h80A571F2;	14'h08FB: data <= 32'h80AC6783;	14'h08FC: data <= 32'h80B381AE;	14'h08FD: data <= 32'h80BAC071;	14'h08FE: data <= 32'h80C223CA;	14'h08FF: data <= 32'h80C9ABB8;	14'h0900: data <= 32'h80D15838;	14'h0901: data <= 32'h80D92947;	14'h0902: data <= 32'h80E11EE4;	14'h0903: data <= 32'h80E9390C;	14'h0904: data <= 32'h80F177BD;	14'h0905: data <= 32'h80F9DAF4;	14'h0906: data <= 32'h810262AF;	14'h0907: data <= 32'h810B0EED;	14'h0908: data <= 32'h8113DFA9;	14'h0909: data <= 32'h811CD4E2;	14'h090A: data <= 32'h8125EE95;	14'h090B: data <= 32'h812F2CBF;	14'h090C: data <= 32'h81388F5E;	14'h090D: data <= 32'h8142166F;	14'h090E: data <= 32'h814BC1EF;	14'h090F: data <= 32'h815591DC;	14'h0910: data <= 32'h815F8633;	14'h0911: data <= 32'h81699EF1;	14'h0912: data <= 32'h8173DC12;	14'h0913: data <= 32'h817E3D95;	14'h0914: data <= 32'h8188C375;	14'h0915: data <= 32'h81936DB1;	14'h0916: data <= 32'h819E3C44;	14'h0917: data <= 32'h81A92F2D;	14'h0918: data <= 32'h81B44667;	14'h0919: data <= 32'h81BF81EF;	14'h091A: data <= 32'h81CAE1C3;	14'h091B: data <= 32'h81D665DF;	14'h091C: data <= 32'h81E20E3F;	14'h091D: data <= 32'h81EDDAE1;	14'h091E: data <= 32'h81F9CBC1;	14'h091F: data <= 32'h8205E0DB;	14'h0920: data <= 32'h82121A2C;	14'h0921: data <= 32'h821E77B1;	14'h0922: data <= 32'h822AF966;	14'h0923: data <= 32'h82379F47;	14'h0924: data <= 32'h82446951;	14'h0925: data <= 32'h82515780;	14'h0926: data <= 32'h825E69D0;	14'h0927: data <= 32'h826BA03E;	14'h0928: data <= 32'h8278FAC6;	14'h0929: data <= 32'h82867963;	14'h092A: data <= 32'h82941C13;	14'h092B: data <= 32'h82A1E2D1;	14'h092C: data <= 32'h82AFCD99;	14'h092D: data <= 32'h82BDDC67;	14'h092E: data <= 32'h82CC0F38;	14'h092F: data <= 32'h82DA6606;	14'h0930: data <= 32'h82E8E0CE;	14'h0931: data <= 32'h82F77F8D;	14'h0932: data <= 32'h8306423C;	14'h0933: data <= 32'h831528D9;	14'h0934: data <= 32'h83243360;	14'h0935: data <= 32'h833361CA;	14'h0936: data <= 32'h8342B416;	14'h0937: data <= 32'h83522A3D;	14'h0938: data <= 32'h8361C43C;	14'h0939: data <= 32'h8371820D;	14'h093A: data <= 32'h838163AD;	14'h093B: data <= 32'h83916918;	14'h093C: data <= 32'h83A19247;	14'h093D: data <= 32'h83B1DF37;	14'h093E: data <= 32'h83C24FE4;	14'h093F: data <= 32'h83D2E447;	14'h0940: data <= 32'h83E39C5D;	14'h0941: data <= 32'h83F47821;	14'h0942: data <= 32'h8405778D;	14'h0943: data <= 32'h84169A9E;	14'h0944: data <= 32'h8427E14D;	14'h0945: data <= 32'h84394B97;	14'h0946: data <= 32'h844AD976;	14'h0947: data <= 32'h845C8AE4;	14'h0948: data <= 32'h846E5FDE;	14'h0949: data <= 32'h8480585D;	14'h094A: data <= 32'h8492745E;	14'h094B: data <= 32'h84A4B3D9;	14'h094C: data <= 32'h84B716CB;	14'h094D: data <= 32'h84C99D2E;	14'h094E: data <= 32'h84DC46FC;	14'h094F: data <= 32'h84EF1430;	14'h0950: data <= 32'h850204C6;	14'h0951: data <= 32'h851518B6;	14'h0952: data <= 32'h85284FFD;	14'h0953: data <= 32'h853BAA94;	14'h0954: data <= 32'h854F2875;	14'h0955: data <= 32'h8562C99C;	14'h0956: data <= 32'h85768E03;	14'h0957: data <= 32'h858A75A3;	14'h0958: data <= 32'h859E8077;	14'h0959: data <= 32'h85B2AE7A;	14'h095A: data <= 32'h85C6FFA6;	14'h095B: data <= 32'h85DB73F4;	14'h095C: data <= 32'h85F00B5F;	14'h095D: data <= 32'h8604C5E1;	14'h095E: data <= 32'h8619A374;	14'h095F: data <= 32'h862EA412;	14'h0960: data <= 32'h8643C7B4;	14'h0961: data <= 32'h86590E56;	14'h0962: data <= 32'h866E77F1;	14'h0963: data <= 32'h8684047E;	14'h0964: data <= 32'h8699B3F7;	14'h0965: data <= 32'h86AF8657;	14'h0966: data <= 32'h86C57B96;	14'h0967: data <= 32'h86DB93B0;	14'h0968: data <= 32'h86F1CE9C;	14'h0969: data <= 32'h87082C55;	14'h096A: data <= 32'h871EACD5;	14'h096B: data <= 32'h87355014;	14'h096C: data <= 32'h874C160D;	14'h096D: data <= 32'h8762FEB9;	14'h096E: data <= 32'h877A0A12;	14'h096F: data <= 32'h8791380F;	14'h0970: data <= 32'h87A888AC;	14'h0971: data <= 32'h87BFFBE2;	14'h0972: data <= 32'h87D791A8;	14'h0973: data <= 32'h87EF49FA;	14'h0974: data <= 32'h880724CF;	14'h0975: data <= 32'h881F2222;	14'h0976: data <= 32'h883741EB;	14'h0977: data <= 32'h884F8423;	14'h0978: data <= 32'h8867E8C4;	14'h0979: data <= 32'h88806FC5;	14'h097A: data <= 32'h88991921;	14'h097B: data <= 32'h88B1E4D1;	14'h097C: data <= 32'h88CAD2CC;	14'h097D: data <= 32'h88E3E30C;	14'h097E: data <= 32'h88FD158A;	14'h097F: data <= 32'h89166A3E;	14'h0980: data <= 32'h892FE121;	14'h0981: data <= 32'h89497A2C;	14'h0982: data <= 32'h89633558;	14'h0983: data <= 32'h897D129C;	14'h0984: data <= 32'h899711F3;	14'h0985: data <= 32'h89B13353;	14'h0986: data <= 32'h89CB76B6;	14'h0987: data <= 32'h89E5DC14;	14'h0988: data <= 32'h8A006366;	14'h0989: data <= 32'h8A1B0CA3;	14'h098A: data <= 32'h8A35D7C5;	14'h098B: data <= 32'h8A50C4C3;	14'h098C: data <= 32'h8A6BD396;	14'h098D: data <= 32'h8A870436;	14'h098E: data <= 32'h8AA2569B;	14'h098F: data <= 32'h8ABDCABD;	14'h0990: data <= 32'h8AD96095;	14'h0991: data <= 32'h8AF5181B;	14'h0992: data <= 32'h8B10F145;	14'h0993: data <= 32'h8B2CEC0E;	14'h0994: data <= 32'h8B49086C;	14'h0995: data <= 32'h8B654657;	14'h0996: data <= 32'h8B81A5C7;	14'h0997: data <= 32'h8B9E26B5;	14'h0998: data <= 32'h8BBAC918;	14'h0999: data <= 32'h8BD78CE7;	14'h099A: data <= 32'h8BF4721B;	14'h099B: data <= 32'h8C1178AA;	14'h099C: data <= 32'h8C2EA08E;	14'h099D: data <= 32'h8C4BE9BD;	14'h099E: data <= 32'h8C69542F;	14'h099F: data <= 32'h8C86DFDB;	14'h09A0: data <= 32'h8CA48CBA;	14'h09A1: data <= 32'h8CC25AC2;	14'h09A2: data <= 32'h8CE049EB;	14'h09A3: data <= 32'h8CFE5A2C;	14'h09A4: data <= 32'h8D1C8B7D;	14'h09A5: data <= 32'h8D3ADDD5;	14'h09A6: data <= 32'h8D59512B;	14'h09A7: data <= 32'h8D77E577;	14'h09A8: data <= 32'h8D969AAF;	14'h09A9: data <= 32'h8DB570CB;	14'h09AA: data <= 32'h8DD467C3;	14'h09AB: data <= 32'h8DF37F8C;	14'h09AC: data <= 32'h8E12B81F;	14'h09AD: data <= 32'h8E321172;	14'h09AE: data <= 32'h8E518B7C;	14'h09AF: data <= 32'h8E712635;	14'h09B0: data <= 32'h8E90E192;	14'h09B1: data <= 32'h8EB0BD8C;	14'h09B2: data <= 32'h8ED0BA18;	14'h09B3: data <= 32'h8EF0D72E;	14'h09B4: data <= 32'h8F1114C4;	14'h09B5: data <= 32'h8F3172D1;	14'h09B6: data <= 32'h8F51F14C;	14'h09B7: data <= 32'h8F72902C;	14'h09B8: data <= 32'h8F934F66;	14'h09B9: data <= 32'h8FB42EF3;	14'h09BA: data <= 32'h8FD52EC7;	14'h09BB: data <= 32'h8FF64EDB;	14'h09BC: data <= 32'h90178F23;	14'h09BD: data <= 32'h9038EF97;	14'h09BE: data <= 32'h905A702D;	14'h09BF: data <= 32'h907C10DC;	14'h09C0: data <= 32'h909DD199;	14'h09C1: data <= 32'h90BFB25C;	14'h09C2: data <= 32'h90E1B31A;	14'h09C3: data <= 32'h9103D3C9;	14'h09C4: data <= 32'h91261460;	14'h09C5: data <= 32'h914874D5;	14'h09C6: data <= 32'h916AF51E;	14'h09C7: data <= 32'h918D9531;	14'h09C8: data <= 32'h91B05504;	14'h09C9: data <= 32'h91D3348D;	14'h09CA: data <= 32'h91F633C3;	14'h09CB: data <= 32'h9219529A;	14'h09CC: data <= 32'h923C9109;	14'h09CD: data <= 32'h925FEF07;	14'h09CE: data <= 32'h92836C88;	14'h09CF: data <= 32'h92A70982;	14'h09D0: data <= 32'h92CAC5EB;	14'h09D1: data <= 32'h92EEA1BA;	14'h09D2: data <= 32'h93129CE3;	14'h09D3: data <= 32'h9336B75D;	14'h09D4: data <= 32'h935AF11C;	14'h09D5: data <= 32'h937F4A17;	14'h09D6: data <= 32'h93A3C243;	14'h09D7: data <= 32'h93C85995;	14'h09D8: data <= 32'h93ED1004;	14'h09D9: data <= 32'h9411E584;	14'h09DA: data <= 32'h9436DA0B;	14'h09DB: data <= 32'h945BED8E;	14'h09DC: data <= 32'h94812003;	14'h09DD: data <= 32'h94A6715F;	14'h09DE: data <= 32'h94CBE197;	14'h09DF: data <= 32'h94F170A0;	14'h09E0: data <= 32'h95171E70;	14'h09E1: data <= 32'h953CEAFC;	14'h09E2: data <= 32'h9562D639;	14'h09E3: data <= 32'h9588E01C;	14'h09E4: data <= 32'h95AF089A;	14'h09E5: data <= 32'h95D54FA8;	14'h09E6: data <= 32'h95FBB53B;	14'h09E7: data <= 32'h96223948;	14'h09E8: data <= 32'h9648DBC5;	14'h09E9: data <= 32'h966F9CA5;	14'h09EA: data <= 32'h96967BDE;	14'h09EB: data <= 32'h96BD7965;	14'h09EC: data <= 32'h96E4952E;	14'h09ED: data <= 32'h970BCF2E;	14'h09EE: data <= 32'h9733275B;	14'h09EF: data <= 32'h975A9DA7;	14'h09F0: data <= 32'h97823209;	14'h09F1: data <= 32'h97A9E475;	14'h09F2: data <= 32'h97D1B4DF;	14'h09F3: data <= 32'h97F9A33C;	14'h09F4: data <= 32'h9821AF81;	14'h09F5: data <= 32'h9849D9A2;	14'h09F6: data <= 32'h98722193;	14'h09F7: data <= 32'h989A8749;	14'h09F8: data <= 32'h98C30AB8;	14'h09F9: data <= 32'h98EBABD5;	14'h09FA: data <= 32'h99146A94;	14'h09FB: data <= 32'h993D46E9;	14'h09FC: data <= 32'h996640C9;	14'h09FD: data <= 32'h998F5827;	14'h09FE: data <= 32'h99B88CF8;	14'h09FF: data <= 32'h99E1DF30;	14'h0A00: data <= 32'h9A0B4EC3;	14'h0A01: data <= 32'h9A34DBA6;	14'h0A02: data <= 32'h9A5E85CC;	14'h0A03: data <= 32'h9A884D29;	14'h0A04: data <= 32'h9AB231B1;	14'h0A05: data <= 32'h9ADC3359;	14'h0A06: data <= 32'h9B065214;	14'h0A07: data <= 32'h9B308DD6;	14'h0A08: data <= 32'h9B5AE693;	14'h0A09: data <= 32'h9B855C3E;	14'h0A0A: data <= 32'h9BAFEECD;	14'h0A0B: data <= 32'h9BDA9E31;	14'h0A0C: data <= 32'h9C056A60;	14'h0A0D: data <= 32'h9C30534C;	14'h0A0E: data <= 32'h9C5B58EA;	14'h0A0F: data <= 32'h9C867B2D;	14'h0A10: data <= 32'h9CB1BA08;	14'h0A11: data <= 32'h9CDD1570;	14'h0A12: data <= 32'h9D088D58;	14'h0A13: data <= 32'h9D3421B2;	14'h0A14: data <= 32'h9D5FD274;	14'h0A15: data <= 32'h9D8B9F8F;	14'h0A16: data <= 32'h9DB788F9;	14'h0A17: data <= 32'h9DE38EA3;	14'h0A18: data <= 32'h9E0FB081;	14'h0A19: data <= 32'h9E3BEE87;	14'h0A1A: data <= 32'h9E6848A8;	14'h0A1B: data <= 32'h9E94BED7;	14'h0A1C: data <= 32'h9EC15108;	14'h0A1D: data <= 32'h9EEDFF2D;	14'h0A1E: data <= 32'h9F1AC93A;	14'h0A1F: data <= 32'h9F47AF21;	14'h0A20: data <= 32'h9F74B0D7;	14'h0A21: data <= 32'h9FA1CE4D;	14'h0A22: data <= 32'h9FCF0778;	14'h0A23: data <= 32'h9FFC5C49;	14'h0A24: data <= 32'hA029CCB4;	14'h0A25: data <= 32'hA05758AD;	14'h0A26: data <= 32'hA0850025;	14'h0A27: data <= 32'hA0B2C310;	14'h0A28: data <= 32'hA0E0A160;	14'h0A29: data <= 32'hA10E9B09;	14'h0A2A: data <= 32'hA13CAFFD;	14'h0A2B: data <= 32'hA16AE02F;	14'h0A2C: data <= 32'hA1992B92;	14'h0A2D: data <= 32'hA1C79217;	14'h0A2E: data <= 32'hA1F613B3;	14'h0A2F: data <= 32'hA224B057;	14'h0A30: data <= 32'hA25367F7;	14'h0A31: data <= 32'hA2823A84;	14'h0A32: data <= 32'hA2B127F2;	14'h0A33: data <= 32'hA2E03032;	14'h0A34: data <= 32'hA30F5338;	14'h0A35: data <= 32'hA33E90F6;	14'h0A36: data <= 32'hA36DE95D;	14'h0A37: data <= 32'hA39D5C62;	14'h0A38: data <= 32'hA3CCE9F5;	14'h0A39: data <= 32'hA3FC9209;	14'h0A3A: data <= 32'hA42C5491;	14'h0A3B: data <= 32'hA45C317F;	14'h0A3C: data <= 32'hA48C28C5;	14'h0A3D: data <= 32'hA4BC3A55;	14'h0A3E: data <= 32'hA4EC6621;	14'h0A3F: data <= 32'hA51CAC1D;	14'h0A40: data <= 32'hA54D0C39;	14'h0A41: data <= 32'hA57D8667;	14'h0A42: data <= 32'hA5AE1A9B;	14'h0A43: data <= 32'hA5DEC8C5;	14'h0A44: data <= 32'hA60F90D9;	14'h0A45: data <= 32'hA64072C7;	14'h0A46: data <= 32'hA6716E82;	14'h0A47: data <= 32'hA6A283FC;	14'h0A48: data <= 32'hA6D3B327;	14'h0A49: data <= 32'hA704FBF4;	14'h0A4A: data <= 32'hA7365E56;	14'h0A4B: data <= 32'hA767DA3D;	14'h0A4C: data <= 32'hA7996F9D;	14'h0A4D: data <= 32'hA7CB1E66;	14'h0A4E: data <= 32'hA7FCE68B;	14'h0A4F: data <= 32'hA82EC7FC;	14'h0A50: data <= 32'hA860C2AD;	14'h0A51: data <= 32'hA892D68E;	14'h0A52: data <= 32'hA8C50391;	14'h0A53: data <= 32'hA8F749A7;	14'h0A54: data <= 32'hA929A8C2;	14'h0A55: data <= 32'hA95C20D5;	14'h0A56: data <= 32'hA98EB1CF;	14'h0A57: data <= 32'hA9C15BA3;	14'h0A58: data <= 32'hA9F41E41;	14'h0A59: data <= 32'hAA26F99D;	14'h0A5A: data <= 32'hAA59EDA6;	14'h0A5B: data <= 32'hAA8CFA4E;	14'h0A5C: data <= 32'hAAC01F86;	14'h0A5D: data <= 32'hAAF35D41;	14'h0A5E: data <= 32'hAB26B36E;	14'h0A5F: data <= 32'hAB5A2200;	14'h0A60: data <= 32'hAB8DA8E7;	14'h0A61: data <= 32'hABC14815;	14'h0A62: data <= 32'hABF4FF7B;	14'h0A63: data <= 32'hAC28CF0A;	14'h0A64: data <= 32'hAC5CB6B3;	14'h0A65: data <= 32'hAC90B667;	14'h0A66: data <= 32'hACC4CE17;	14'h0A67: data <= 32'hACF8FDB5;	14'h0A68: data <= 32'hAD2D4530;	14'h0A69: data <= 32'hAD61A47B;	14'h0A6A: data <= 32'hAD961B86;	14'h0A6B: data <= 32'hADCAAA43;	14'h0A6C: data <= 32'hADFF50A1;	14'h0A6D: data <= 32'hAE340E92;	14'h0A6E: data <= 32'hAE68E406;	14'h0A6F: data <= 32'hAE9DD0EF;	14'h0A70: data <= 32'hAED2D53E;	14'h0A71: data <= 32'hAF07F0E2;	14'h0A72: data <= 32'hAF3D23CD;	14'h0A73: data <= 32'hAF726DF0;	14'h0A74: data <= 32'hAFA7CF3B;	14'h0A75: data <= 32'hAFDD479E;	14'h0A76: data <= 32'hB012D70B;	14'h0A77: data <= 32'hB0487D72;	14'h0A78: data <= 32'hB07E3AC4;	14'h0A79: data <= 32'hB0B40EF1;	14'h0A7A: data <= 32'hB0E9F9E9;	14'h0A7B: data <= 32'hB11FFB9E;	14'h0A7C: data <= 32'hB15613FF;	14'h0A7D: data <= 32'hB18C42FE;	14'h0A7E: data <= 32'hB1C2888A;	14'h0A7F: data <= 32'hB1F8E493;	14'h0A80: data <= 32'hB22F570C;	14'h0A81: data <= 32'hB265DFE3;	14'h0A82: data <= 32'hB29C7F08;	14'h0A83: data <= 32'hB2D3346D;	14'h0A84: data <= 32'hB30A0002;	14'h0A85: data <= 32'hB340E1B6;	14'h0A86: data <= 32'hB377D97B;	14'h0A87: data <= 32'hB3AEE740;	14'h0A88: data <= 32'hB3E60AF5;	14'h0A89: data <= 32'hB41D448A;	14'h0A8A: data <= 32'hB45493F0;	14'h0A8B: data <= 32'hB48BF917;	14'h0A8C: data <= 32'hB4C373EF;	14'h0A8D: data <= 32'hB4FB0468;	14'h0A8E: data <= 32'hB532AA72;	14'h0A8F: data <= 32'hB56A65FC;	14'h0A90: data <= 32'hB5A236F8;	14'h0A91: data <= 32'hB5DA1D54;	14'h0A92: data <= 32'hB6121901;	14'h0A93: data <= 32'hB64A29EF;	14'h0A94: data <= 32'hB682500D;	14'h0A95: data <= 32'hB6BA8B4C;	14'h0A96: data <= 32'hB6F2DB9B;	14'h0A97: data <= 32'hB72B40EA;	14'h0A98: data <= 32'hB763BB29;	14'h0A99: data <= 32'hB79C4A47;	14'h0A9A: data <= 32'hB7D4EE35;	14'h0A9B: data <= 32'hB80DA6E2;	14'h0A9C: data <= 32'hB846743E;	14'h0A9D: data <= 32'hB87F5638;	14'h0A9E: data <= 32'hB8B84CC1;	14'h0A9F: data <= 32'hB8F157C7;	14'h0AA0: data <= 32'hB92A773A;	14'h0AA1: data <= 32'hB963AB0A;	14'h0AA2: data <= 32'hB99CF327;	14'h0AA3: data <= 32'hB9D64F80;	14'h0AA4: data <= 32'hBA0FC004;	14'h0AA5: data <= 32'hBA4944A3;	14'h0AA6: data <= 32'hBA82DD4D;	14'h0AA7: data <= 32'hBABC89F1;	14'h0AA8: data <= 32'hBAF64A7D;	14'h0AA9: data <= 32'hBB301EE3;	14'h0AAA: data <= 32'hBB6A0711;	14'h0AAB: data <= 32'hBBA402F6;	14'h0AAC: data <= 32'hBBDE1282;	14'h0AAD: data <= 32'hBC1835A4;	14'h0AAE: data <= 32'hBC526C4B;	14'h0AAF: data <= 32'hBC8CB667;	14'h0AB0: data <= 32'hBCC713E7;	14'h0AB1: data <= 32'hBD0184BA;	14'h0AB2: data <= 32'hBD3C08CF;	14'h0AB3: data <= 32'hBD76A016;	14'h0AB4: data <= 32'hBDB14A7D;	14'h0AB5: data <= 32'hBDEC07F4;	14'h0AB6: data <= 32'hBE26D86A;	14'h0AB7: data <= 32'hBE61BBCE;	14'h0AB8: data <= 32'hBE9CB20F;	14'h0AB9: data <= 32'hBED7BB1D;	14'h0ABA: data <= 32'hBF12D6E5;	14'h0ABB: data <= 32'hBF4E0557;	14'h0ABC: data <= 32'hBF894663;	14'h0ABD: data <= 32'hBFC499F6;	14'h0ABE: data <= 32'hC0000001;	14'h0ABF: data <= 32'hC03B7872;	14'h0AC0: data <= 32'hC0770337;	14'h0AC1: data <= 32'hC0B2A040;	14'h0AC2: data <= 32'hC0EE4F7C;	14'h0AC3: data <= 32'hC12A10D9;	14'h0AC4: data <= 32'hC165E447;	14'h0AC5: data <= 32'hC1A1C9B4;	14'h0AC6: data <= 32'hC1DDC10E;	14'h0AC7: data <= 32'hC219CA45;	14'h0AC8: data <= 32'hC255E547;	14'h0AC9: data <= 32'hC2921204;	14'h0ACA: data <= 32'hC2CE5069;	14'h0ACB: data <= 32'hC30AA066;	14'h0ACC: data <= 32'hC34701E9;	14'h0ACD: data <= 32'hC38374E1;	14'h0ACE: data <= 32'hC3BFF93C;	14'h0ACF: data <= 32'hC3FC8EE9;	14'h0AD0: data <= 32'hC43935D6;	14'h0AD1: data <= 32'hC475EDF3;	14'h0AD2: data <= 32'hC4B2B72D;	14'h0AD3: data <= 32'hC4EF9174;	14'h0AD4: data <= 32'hC52C7CB5;	14'h0AD5: data <= 32'hC56978E0;	14'h0AD6: data <= 32'hC5A685E2;	14'h0AD7: data <= 32'hC5E3A3AA;	14'h0AD8: data <= 32'hC620D227;	14'h0AD9: data <= 32'hC65E1147;	14'h0ADA: data <= 32'hC69B60F8;	14'h0ADB: data <= 32'hC6D8C129;	14'h0ADC: data <= 32'hC71631C8;	14'h0ADD: data <= 32'hC753B2C4;	14'h0ADE: data <= 32'hC791440A;	14'h0ADF: data <= 32'hC7CEE589;	14'h0AE0: data <= 32'hC80C9730;	14'h0AE1: data <= 32'hC84A58EC;	14'h0AE2: data <= 32'hC8882AAC;	14'h0AE3: data <= 32'hC8C60C5E;	14'h0AE4: data <= 32'hC903FDF0;	14'h0AE5: data <= 32'hC941FF51;	14'h0AE6: data <= 32'hC980106F;	14'h0AE7: data <= 32'hC9BE3137;	14'h0AE8: data <= 32'hC9FC6198;	14'h0AE9: data <= 32'hCA3AA180;	14'h0AEA: data <= 32'hCA78F0DE;	14'h0AEB: data <= 32'hCAB74F9F;	14'h0AEC: data <= 32'hCAF5BDB1;	14'h0AED: data <= 32'hCB343B02;	14'h0AEE: data <= 32'hCB72C781;	14'h0AEF: data <= 32'hCBB1631B;	14'h0AF0: data <= 32'hCBF00DBF;	14'h0AF1: data <= 32'hCC2EC75A;	14'h0AF2: data <= 32'hCC6D8FDB;	14'h0AF3: data <= 32'hCCAC672E;	14'h0AF4: data <= 32'hCCEB4D44;	14'h0AF5: data <= 32'hCD2A4208;	14'h0AF6: data <= 32'hCD694569;	14'h0AF7: data <= 32'hCDA85756;	14'h0AF8: data <= 32'hCDE777BB;	14'h0AF9: data <= 32'hCE26A687;	14'h0AFA: data <= 32'hCE65E3A8;	14'h0AFB: data <= 32'hCEA52F0B;	14'h0AFC: data <= 32'hCEE4889E;	14'h0AFD: data <= 32'hCF23F04F;	14'h0AFE: data <= 32'hCF63660B;	14'h0AFF: data <= 32'hCFA2E9C2;	14'h0B00: data <= 32'hCFE27B5F;	14'h0B01: data <= 32'hD0221AD2;	14'h0B02: data <= 32'hD061C807;	14'h0B03: data <= 32'hD0A182EC;	14'h0B04: data <= 32'hD0E14B70;	14'h0B05: data <= 32'hD121217F;	14'h0B06: data <= 32'hD1610507;	14'h0B07: data <= 32'hD1A0F5F7;	14'h0B08: data <= 32'hD1E0F43B;	14'h0B09: data <= 32'hD220FFC1;	14'h0B0A: data <= 32'hD2611877;	14'h0B0B: data <= 32'hD2A13E4B;	14'h0B0C: data <= 32'hD2E17129;	14'h0B0D: data <= 32'hD321B100;	14'h0B0E: data <= 32'hD361FDBD;	14'h0B0F: data <= 32'hD3A2574D;	14'h0B10: data <= 32'hD3E2BD9F;	14'h0B11: data <= 32'hD423309F;	14'h0B12: data <= 32'hD463B03B;	14'h0B13: data <= 32'hD4A43C60;	14'h0B14: data <= 32'hD4E4D4FC;	14'h0B15: data <= 32'hD52579FD;	14'h0B16: data <= 32'hD5662B4F;	14'h0B17: data <= 32'hD5A6E8E1;	14'h0B18: data <= 32'hD5E7B29F;	14'h0B19: data <= 32'hD6288876;	14'h0B1A: data <= 32'hD6696A56;	14'h0B1B: data <= 32'hD6AA5829;	14'h0B1C: data <= 32'hD6EB51DF;	14'h0B1D: data <= 32'hD72C5764;	14'h0B1E: data <= 32'hD76D68A5;	14'h0B1F: data <= 32'hD7AE8591;	14'h0B20: data <= 32'hD7EFAE13;	14'h0B21: data <= 32'hD830E21A;	14'h0B22: data <= 32'hD8722192;	14'h0B23: data <= 32'hD8B36C6A;	14'h0B24: data <= 32'hD8F4C28E;	14'h0B25: data <= 32'hD93623EA;	14'h0B26: data <= 32'hD977906E;	14'h0B27: data <= 32'hD9B90805;	14'h0B28: data <= 32'hD9FA8A9E;	14'h0B29: data <= 32'hDA3C1824;	14'h0B2A: data <= 32'hDA7DB086;	14'h0B2B: data <= 32'hDABF53B0;	14'h0B2C: data <= 32'hDB01018F;	14'h0B2D: data <= 32'hDB42BA11;	14'h0B2E: data <= 32'hDB847D23;	14'h0B2F: data <= 32'hDBC64AB2;	14'h0B30: data <= 32'hDC0822AB;	14'h0B31: data <= 32'hDC4A04FB;	14'h0B32: data <= 32'hDC8BF18E;	14'h0B33: data <= 32'hDCCDE853;	14'h0B34: data <= 32'hDD0FE937;	14'h0B35: data <= 32'hDD51F425;	14'h0B36: data <= 32'hDD94090B;	14'h0B37: data <= 32'hDDD627D7;	14'h0B38: data <= 32'hDE185075;	14'h0B39: data <= 32'hDE5A82D2;	14'h0B3A: data <= 32'hDE9CBEDB;	14'h0B3B: data <= 32'hDEDF047E;	14'h0B3C: data <= 32'hDF2153A6;	14'h0B3D: data <= 32'hDF63AC41;	14'h0B3E: data <= 32'hDFA60E3D;	14'h0B3F: data <= 32'hDFE87985;	14'h0B40: data <= 32'hE02AEE07;	14'h0B41: data <= 32'hE06D6BAF;	14'h0B42: data <= 32'hE0AFF26B;	14'h0B43: data <= 32'hE0F28228;	14'h0B44: data <= 32'hE1351AD1;	14'h0B45: data <= 32'hE177BC55;	14'h0B46: data <= 32'hE1BA66A0;	14'h0B47: data <= 32'hE1FD199E;	14'h0B48: data <= 32'hE23FD53E;	14'h0B49: data <= 32'hE282996A;	14'h0B4A: data <= 32'hE2C56611;	14'h0B4B: data <= 32'hE3083B1F;	14'h0B4C: data <= 32'hE34B1881;	14'h0B4D: data <= 32'hE38DFE23;	14'h0B4E: data <= 32'hE3D0EBF3;	14'h0B4F: data <= 32'hE413E1DD;	14'h0B50: data <= 32'hE456DFCE;	14'h0B51: data <= 32'hE499E5B2;	14'h0B52: data <= 32'hE4DCF377;	14'h0B53: data <= 32'hE5200909;	14'h0B54: data <= 32'hE5632654;	14'h0B55: data <= 32'hE5A64B47;	14'h0B56: data <= 32'hE5E977CC;	14'h0B57: data <= 32'hE62CABD1;	14'h0B58: data <= 32'hE66FE743;	14'h0B59: data <= 32'hE6B32A0E;	14'h0B5A: data <= 32'hE6F6741F;	14'h0B5B: data <= 32'hE739C563;	14'h0B5C: data <= 32'hE77D1DC6;	14'h0B5D: data <= 32'hE7C07D34;	14'h0B5E: data <= 32'hE803E39C;	14'h0B5F: data <= 32'hE84750E8;	14'h0B60: data <= 32'hE88AC506;	14'h0B61: data <= 32'hE8CE3FE2;	14'h0B62: data <= 32'hE911C16A;	14'h0B63: data <= 32'hE9554989;	14'h0B64: data <= 32'hE998D82C;	14'h0B65: data <= 32'hE9DC6D3F;	14'h0B66: data <= 32'hEA2008B0;	14'h0B67: data <= 32'hEA63AA6B;	14'h0B68: data <= 32'hEAA7525C;	14'h0B69: data <= 32'hEAEB0070;	14'h0B6A: data <= 32'hEB2EB494;	14'h0B6B: data <= 32'hEB726EB3;	14'h0B6C: data <= 32'hEBB62EBC;	14'h0B6D: data <= 32'hEBF9F499;	14'h0B6E: data <= 32'hEC3DC038;	14'h0B6F: data <= 32'hEC819185;	14'h0B70: data <= 32'hECC5686D;	14'h0B71: data <= 32'hED0944DB;	14'h0B72: data <= 32'hED4D26BE;	14'h0B73: data <= 32'hED910E00;	14'h0B74: data <= 32'hEDD4FA8F;	14'h0B75: data <= 32'hEE18EC57;	14'h0B76: data <= 32'hEE5CE345;	14'h0B77: data <= 32'hEEA0DF44;	14'h0B78: data <= 32'hEEE4E042;	14'h0B79: data <= 32'hEF28E62B;	14'h0B7A: data <= 32'hEF6CF0EB;	14'h0B7B: data <= 32'hEFB1006F;	14'h0B7C: data <= 32'hEFF514A3;	14'h0B7D: data <= 32'hF0392D74;	14'h0B7E: data <= 32'hF07D4ACE;	14'h0B7F: data <= 32'hF0C16C9D;	14'h0B80: data <= 32'hF10592CE;	14'h0B81: data <= 32'hF149BD4D;	14'h0B82: data <= 32'hF18DEC08;	14'h0B83: data <= 32'hF1D21EE9;	14'h0B84: data <= 32'hF21655DD;	14'h0B85: data <= 32'hF25A90D2;	14'h0B86: data <= 32'hF29ECFB3;	14'h0B87: data <= 32'hF2E3126D;	14'h0B88: data <= 32'hF32758EB;	14'h0B89: data <= 32'hF36BA31B;	14'h0B8A: data <= 32'hF3AFF0E9;	14'h0B8B: data <= 32'hF3F44241;	14'h0B8C: data <= 32'hF438970F;	14'h0B8D: data <= 32'hF47CEF40;	14'h0B8E: data <= 32'hF4C14AC1;	14'h0B8F: data <= 32'hF505A97C;	14'h0B90: data <= 32'hF54A0B60;	14'h0B91: data <= 32'hF58E7058;	14'h0B92: data <= 32'hF5D2D851;	14'h0B93: data <= 32'hF6174337;	14'h0B94: data <= 32'hF65BB0F5;	14'h0B95: data <= 32'hF6A0217A;	14'h0B96: data <= 32'hF6E494B0;	14'h0B97: data <= 32'hF7290A85;	14'h0B98: data <= 32'hF76D82E4;	14'h0B99: data <= 32'hF7B1FDBA;	14'h0B9A: data <= 32'hF7F67AF3;	14'h0B9B: data <= 32'hF83AFA7B;	14'h0B9C: data <= 32'hF87F7C40;	14'h0B9D: data <= 32'hF8C4002C;	14'h0B9E: data <= 32'hF908862D;	14'h0B9F: data <= 32'hF94D0E2E;	14'h0BA0: data <= 32'hF991981D;	14'h0BA1: data <= 32'hF9D623E5;	14'h0BA2: data <= 32'hFA1AB172;	14'h0BA3: data <= 32'hFA5F40B1;	14'h0BA4: data <= 32'hFAA3D18F;	14'h0BA5: data <= 32'hFAE863F7;	14'h0BA6: data <= 32'hFB2CF7D6;	14'h0BA7: data <= 32'hFB718D17;	14'h0BA8: data <= 32'hFBB623A8;	14'h0BA9: data <= 32'hFBFABB75;	14'h0BAA: data <= 32'hFC3F546A;	14'h0BAB: data <= 32'hFC83EE72;	14'h0BAC: data <= 32'hFCC8897B;	14'h0BAD: data <= 32'hFD0D2571;	14'h0BAE: data <= 32'hFD51C240;	14'h0BAF: data <= 32'hFD965FD4;	14'h0BB0: data <= 32'hFDDAFE1A;	14'h0BB1: data <= 32'hFE1F9CFE;	14'h0BB2: data <= 32'hFE643C6B;	14'h0BB3: data <= 32'hFEA8DC4F;	14'h0BB4: data <= 32'hFEED7C96;	14'h0BB5: data <= 32'hFF321D2C;	14'h0BB6: data <= 32'hFF76BDFC;	14'h0BB7: data <= 32'hFFBB5EF5;	14'h0BB8: data <= 32'h00887CBF;	14'h0BB9: data <= 32'h004B8DB2;	14'h0BBA: data <= 32'h000E9EA6;	14'h0BBB: data <= 32'hFFD1AF9B;	14'h0BBC: data <= 32'hFF94C08F;	14'h0BBD: data <= 32'hFF57D183;	14'h0BBE: data <= 32'hFF1AE277;	14'h0BBF: data <= 32'hFEDDF36B;	14'h0BC0: data <= 32'hFEA1045F;	14'h0BC1: data <= 32'hFE641553;	14'h0BC2: data <= 32'hFE272647;	14'h0BC3: data <= 32'hFDEA373B;	14'h0BC4: data <= 32'hFDAD482F;	14'h0BC5: data <= 32'hFD705923;	14'h0BC6: data <= 32'hFD336A17;	14'h0BC7: data <= 32'hFCF67B0A;	14'h0BC8: data <= 32'hFCB98BFE;	14'h0BC9: data <= 32'hFC7C9CF2;	14'h0BCA: data <= 32'hFC3FADE6;	14'h0BCB: data <= 32'hFC02BEDA;	14'h0BCC: data <= 32'hFBC5CFCE;	14'h0BCD: data <= 32'hFB88E0C2;	14'h0BCE: data <= 32'hFB4BF1B6;	14'h0BCF: data <= 32'hFB0F02AA;	14'h0BD0: data <= 32'hFAD2139E;	14'h0BD1: data <= 32'hFA952492;	14'h0BD2: data <= 32'hFA583586;	14'h0BD3: data <= 32'hFA1B467A;	14'h0BD4: data <= 32'hF9DE576E;	14'h0BD5: data <= 32'hF9A16861;	14'h0BD6: data <= 32'hF9647955;	14'h0BD7: data <= 32'hF929E31A;	14'h0BD8: data <= 32'hF8F05218;	14'h0BD9: data <= 32'hF8B6C115;	14'h0BDA: data <= 32'hF87D3013;	14'h0BDB: data <= 32'hF8439F11;	14'h0BDC: data <= 32'hF80A0E0E;	14'h0BDD: data <= 32'hF7D07D0C;	14'h0BDE: data <= 32'hF796EC0A;	14'h0BDF: data <= 32'hF75D5B07;	14'h0BE0: data <= 32'hF723CA05;	14'h0BE1: data <= 32'hF6EA3903;	14'h0BE2: data <= 32'hF6B0A800;	14'h0BE3: data <= 32'hF67716FE;	14'h0BE4: data <= 32'hF63D85FC;	14'h0BE5: data <= 32'hF603F4F9;	14'h0BE6: data <= 32'hF5CA63F7;	14'h0BE7: data <= 32'hF590D2F5;	14'h0BE8: data <= 32'hF55741F3;	14'h0BE9: data <= 32'hF51DB0F0;	14'h0BEA: data <= 32'hF4E41FEE;	14'h0BEB: data <= 32'hF4AA8EEC;	14'h0BEC: data <= 32'hF470FDE9;	14'h0BED: data <= 32'hF4376CE7;	14'h0BEE: data <= 32'hF3FDDBE5;	14'h0BEF: data <= 32'hF3C44AE2;	14'h0BF0: data <= 32'hF38AB9E0;	14'h0BF1: data <= 32'hF35128DE;	14'h0BF2: data <= 32'hF31797DB;	14'h0BF3: data <= 32'hF2DE06D9;	14'h0BF4: data <= 32'hF2A475D7;	14'h0BF5: data <= 32'hF26D3BFB;	14'h0BF6: data <= 32'hF2399BE4;	14'h0BF7: data <= 32'hF205FBCE;	14'h0BF8: data <= 32'hF1D25BB7;	14'h0BF9: data <= 32'hF19EBBA1;	14'h0BFA: data <= 32'hF16B1B8A;	14'h0BFB: data <= 32'hF1377B73;	14'h0BFC: data <= 32'hF103DB5D;	14'h0BFD: data <= 32'hF0D03B46;	14'h0BFE: data <= 32'hF09C9B30;	14'h0BFF: data <= 32'hF068FB19;	14'h0C00: data <= 32'hF0355B02;	14'h0C01: data <= 32'hF001BAEC;	14'h0C02: data <= 32'hEFCE1AD5;	14'h0C03: data <= 32'hEF9A7ABF;	14'h0C04: data <= 32'hEF66DAA8;	14'h0C05: data <= 32'hEF333A91;	14'h0C06: data <= 32'hEEFF9A7B;	14'h0C07: data <= 32'hEECBFA64;	14'h0C08: data <= 32'hEE985A4E;	14'h0C09: data <= 32'hEE64BA37;	14'h0C0A: data <= 32'hEE311A20;	14'h0C0B: data <= 32'hEDFD7A0A;	14'h0C0C: data <= 32'hEDC9D9F3;	14'h0C0D: data <= 32'hED9639DD;	14'h0C0E: data <= 32'hED6299C6;	14'h0C0F: data <= 32'hED2EF9AF;	14'h0C10: data <= 32'hECFB5999;	14'h0C11: data <= 32'hECC7B982;	14'h0C12: data <= 32'hEC94196C;	14'h0C13: data <= 32'hEC613882;	14'h0C14: data <= 32'hEC35CF5B;	14'h0C15: data <= 32'hEC0A6633;	14'h0C16: data <= 32'hEBDEFD0C;	14'h0C17: data <= 32'hEBB393E4;	14'h0C18: data <= 32'hEB882ABC;	14'h0C19: data <= 32'hEB5CC195;	14'h0C1A: data <= 32'hEB31586D;	14'h0C1B: data <= 32'hEB05EF46;	14'h0C1C: data <= 32'hEADA861E;	14'h0C1D: data <= 32'hEAAF1CF7;	14'h0C1E: data <= 32'hEA83B3CF;	14'h0C1F: data <= 32'hEA584AA8;	14'h0C20: data <= 32'hEA2CE180;	14'h0C21: data <= 32'hEA017859;	14'h0C22: data <= 32'hE9D60F31;	14'h0C23: data <= 32'hE9AAA60A;	14'h0C24: data <= 32'hE97F3CE2;	14'h0C25: data <= 32'hE953D3BB;	14'h0C26: data <= 32'hE9286A93;	14'h0C27: data <= 32'hE8FD016C;	14'h0C28: data <= 32'hE8D19844;	14'h0C29: data <= 32'hE8A62F1D;	14'h0C2A: data <= 32'hE87AC5F5;	14'h0C2B: data <= 32'hE84F5CCE;	14'h0C2C: data <= 32'hE823F3A6;	14'h0C2D: data <= 32'hE7F88A7F;	14'h0C2E: data <= 32'hE7CD2157;	14'h0C2F: data <= 32'hE7A1B830;	14'h0C30: data <= 32'hE7764F08;	14'h0C31: data <= 32'hE74AE5E0;	14'h0C32: data <= 32'hE726A6F2;	14'h0C33: data <= 32'hE70455D8;	14'h0C34: data <= 32'hE6E204BE;	14'h0C35: data <= 32'hE6BFB3A3;	14'h0C36: data <= 32'hE69D6289;	14'h0C37: data <= 32'hE67B116F;	14'h0C38: data <= 32'hE658C055;	14'h0C39: data <= 32'hE6366F3B;	14'h0C3A: data <= 32'hE6141E20;	14'h0C3B: data <= 32'hE5F1CD06;	14'h0C3C: data <= 32'hE5CF7BEC;	14'h0C3D: data <= 32'hE5AD2AD2;	14'h0C3E: data <= 32'hE58AD9B8;	14'h0C3F: data <= 32'hE568889D;	14'h0C40: data <= 32'hE5463783;	14'h0C41: data <= 32'hE523E669;	14'h0C42: data <= 32'hE501954F;	14'h0C43: data <= 32'hE4DF4435;	14'h0C44: data <= 32'hE4BCF31A;	14'h0C45: data <= 32'hE49AA200;	14'h0C46: data <= 32'hE47850E6;	14'h0C47: data <= 32'hE455FFCC;	14'h0C48: data <= 32'hE433AEB2;	14'h0C49: data <= 32'hE4115D97;	14'h0C4A: data <= 32'hE3EF0C7D;	14'h0C4B: data <= 32'hE3CCBB63;	14'h0C4C: data <= 32'hE3AA6A49;	14'h0C4D: data <= 32'hE388192F;	14'h0C4E: data <= 32'hE365C814;	14'h0C4F: data <= 32'hE34376FA;	14'h0C50: data <= 32'hE324C44E;	14'h0C51: data <= 32'hE309E9F6;	14'h0C52: data <= 32'hE2EF0F9E;	14'h0C53: data <= 32'hE2D43547;	14'h0C54: data <= 32'hE2B95AEF;	14'h0C55: data <= 32'hE29E8097;	14'h0C56: data <= 32'hE283A640;	14'h0C57: data <= 32'hE268CBE8;	14'h0C58: data <= 32'hE24DF190;	14'h0C59: data <= 32'hE2331739;	14'h0C5A: data <= 32'hE2183CE1;	14'h0C5B: data <= 32'hE1FD6289;	14'h0C5C: data <= 32'hE1E28832;	14'h0C5D: data <= 32'hE1C7ADDA;	14'h0C5E: data <= 32'hE1ACD382;	14'h0C5F: data <= 32'hE191F92A;	14'h0C60: data <= 32'hE1771ED3;	14'h0C61: data <= 32'hE15C447B;	14'h0C62: data <= 32'hE1416A23;	14'h0C63: data <= 32'hE1268FCC;	14'h0C64: data <= 32'hE10BB574;	14'h0C65: data <= 32'hE0F0DB1C;	14'h0C66: data <= 32'hE0D600C5;	14'h0C67: data <= 32'hE0BB266D;	14'h0C68: data <= 32'hE0A04C15;	14'h0C69: data <= 32'hE08571BE;	14'h0C6A: data <= 32'hE06A9766;	14'h0C6B: data <= 32'hE04FBD0E;	14'h0C6C: data <= 32'hE034E2B6;	14'h0C6D: data <= 32'hE01A085F;	14'h0C6E: data <= 32'hDFFFF5B0;	14'h0C6F: data <= 32'hDFE9657C;	14'h0C70: data <= 32'hDFD2D548;	14'h0C71: data <= 32'hDFBC4513;	14'h0C72: data <= 32'hDFA5B4DF;	14'h0C73: data <= 32'hDF8F24AA;	14'h0C74: data <= 32'hDF789476;	14'h0C75: data <= 32'hDF620441;	14'h0C76: data <= 32'hDF4B740D;	14'h0C77: data <= 32'hDF34E3D9;	14'h0C78: data <= 32'hDF1E53A4;	14'h0C79: data <= 32'hDF07C370;	14'h0C7A: data <= 32'hDEF1333B;	14'h0C7B: data <= 32'hDEDAA307;	14'h0C7C: data <= 32'hDEC412D3;	14'h0C7D: data <= 32'hDEAD829E;	14'h0C7E: data <= 32'hDE96F26A;	14'h0C7F: data <= 32'hDE806235;	14'h0C80: data <= 32'hDE69D201;	14'h0C81: data <= 32'hDE5341CC;	14'h0C82: data <= 32'hDE3CB198;	14'h0C83: data <= 32'hDE262164;	14'h0C84: data <= 32'hDE0F912F;	14'h0C85: data <= 32'hDDF900FB;	14'h0C86: data <= 32'hDDE270C6;	14'h0C87: data <= 32'hDDCBE092;	14'h0C88: data <= 32'hDDB5505E;	14'h0C89: data <= 32'hDD9EC029;	14'h0C8A: data <= 32'hDD882FF5;	14'h0C8B: data <= 32'hDD719FC0;	14'h0C8C: data <= 32'hDD5B0F8C;	14'h0C8D: data <= 32'hDD44FCCC;	14'h0C8E: data <= 32'hDD2EFB59;	14'h0C8F: data <= 32'hDD18F9E7;	14'h0C90: data <= 32'hDD02F874;	14'h0C91: data <= 32'hDCECF702;	14'h0C92: data <= 32'hDCD6F590;	14'h0C93: data <= 32'hDCC0F41D;	14'h0C94: data <= 32'hDCAAF2AB;	14'h0C95: data <= 32'hDC94F138;	14'h0C96: data <= 32'hDC7EEFC6;	14'h0C97: data <= 32'hDC68EE54;	14'h0C98: data <= 32'hDC52ECE1;	14'h0C99: data <= 32'hDC3CEB6F;	14'h0C9A: data <= 32'hDC26E9FC;	14'h0C9B: data <= 32'hDC10E88A;	14'h0C9C: data <= 32'hDBFAE718;	14'h0C9D: data <= 32'hDBE4E5A5;	14'h0C9E: data <= 32'hDBCEE433;	14'h0C9F: data <= 32'hDBB8E2C0;	14'h0CA0: data <= 32'hDBA2E14E;	14'h0CA1: data <= 32'hDB8CDFDC;	14'h0CA2: data <= 32'hDB76DE69;	14'h0CA3: data <= 32'hDB60DCF7;	14'h0CA4: data <= 32'hDB4ADB84;	14'h0CA5: data <= 32'hDB34DA12;	14'h0CA6: data <= 32'hDB1ED8A0;	14'h0CA7: data <= 32'hDB08D72D;	14'h0CA8: data <= 32'hDAF2D5BB;	14'h0CA9: data <= 32'hDADCD448;	14'h0CAA: data <= 32'hDAC6D2D6;	14'h0CAB: data <= 32'hDAAF3342;	14'h0CAC: data <= 32'hDA966288;	14'h0CAD: data <= 32'hDA7D91CE;	14'h0CAE: data <= 32'hDA64C114;	14'h0CAF: data <= 32'hDA4BF05A;	14'h0CB0: data <= 32'hDA331F9F;	14'h0CB1: data <= 32'hDA1A4EE5;	14'h0CB2: data <= 32'hDA017E2B;	14'h0CB3: data <= 32'hD9E8AD71;	14'h0CB4: data <= 32'hD9CFDCB7;	14'h0CB5: data <= 32'hD9B70BFD;	14'h0CB6: data <= 32'hD99E3B43;	14'h0CB7: data <= 32'hD9856A89;	14'h0CB8: data <= 32'hD96C99CF;	14'h0CB9: data <= 32'hD953C914;	14'h0CBA: data <= 32'hD93AF85A;	14'h0CBB: data <= 32'hD92227A0;	14'h0CBC: data <= 32'hD90956E6;	14'h0CBD: data <= 32'hD8F0862C;	14'h0CBE: data <= 32'hD8D7B572;	14'h0CBF: data <= 32'hD8BEE4B8;	14'h0CC0: data <= 32'hD8A613FE;	14'h0CC1: data <= 32'hD88D4344;	14'h0CC2: data <= 32'hD8747289;	14'h0CC3: data <= 32'hD85BA1CF;	14'h0CC4: data <= 32'hD842D115;	14'h0CC5: data <= 32'hD82A005B;	14'h0CC6: data <= 32'hD8112FA1;	14'h0CC7: data <= 32'hD7F85EE7;	14'h0CC8: data <= 32'hD7DF8E2D;	14'h0CC9: data <= 32'hD7C54297;	14'h0CCA: data <= 32'hD7A704B8;	14'h0CCB: data <= 32'hD788C6D9;	14'h0CCC: data <= 32'hD76A88FA;	14'h0CCD: data <= 32'hD74C4B1B;	14'h0CCE: data <= 32'hD72E0D3C;	14'h0CCF: data <= 32'hD70FCF5D;	14'h0CD0: data <= 32'hD6F1917E;	14'h0CD1: data <= 32'hD6D3539E;	14'h0CD2: data <= 32'hD6B515BF;	14'h0CD3: data <= 32'hD696D7E0;	14'h0CD4: data <= 32'hD6789A01;	14'h0CD5: data <= 32'hD65A5C22;	14'h0CD6: data <= 32'hD63C1E43;	14'h0CD7: data <= 32'hD61DE064;	14'h0CD8: data <= 32'hD5FFA285;	14'h0CD9: data <= 32'hD5E164A6;	14'h0CDA: data <= 32'hD5C326C7;	14'h0CDB: data <= 32'hD5A4E8E8;	14'h0CDC: data <= 32'hD586AB09;	14'h0CDD: data <= 32'hD5686D29;	14'h0CDE: data <= 32'hD54A2F4A;	14'h0CDF: data <= 32'hD52BF16B;	14'h0CE0: data <= 32'hD50DB38C;	14'h0CE1: data <= 32'hD4EF75AD;	14'h0CE2: data <= 32'hD4D137CE;	14'h0CE3: data <= 32'hD4B2F9EF;	14'h0CE4: data <= 32'hD494BC10;	14'h0CE5: data <= 32'hD4767E31;	14'h0CE6: data <= 32'hD4584052;	14'h0CE7: data <= 32'hD43A0273;	14'h0CE8: data <= 32'hD4154765;	14'h0CE9: data <= 32'hD3F0586D;	14'h0CEA: data <= 32'hD3CB6976;	14'h0CEB: data <= 32'hD3A67A7F;	14'h0CEC: data <= 32'hD3818B87;	14'h0CED: data <= 32'hD35C9C90;	14'h0CEE: data <= 32'hD337AD98;	14'h0CEF: data <= 32'hD312BEA1;	14'h0CF0: data <= 32'hD2EDCFAA;	14'h0CF1: data <= 32'hD2C8E0B2;	14'h0CF2: data <= 32'hD2A3F1BB;	14'h0CF3: data <= 32'hD27F02C3;	14'h0CF4: data <= 32'hD25A13CC;	14'h0CF5: data <= 32'hD23524D5;	14'h0CF6: data <= 32'hD21035DD;	14'h0CF7: data <= 32'hD1EB46E6;	14'h0CF8: data <= 32'hD1C657EE;	14'h0CF9: data <= 32'hD1A168F7;	14'h0CFA: data <= 32'hD17C7A00;	14'h0CFB: data <= 32'hD1578B08;	14'h0CFC: data <= 32'hD1329C11;	14'h0CFD: data <= 32'hD10DAD19;	14'h0CFE: data <= 32'hD0E8BE22;	14'h0CFF: data <= 32'hD0C3CF2B;	14'h0D00: data <= 32'hD09EE033;	14'h0D01: data <= 32'hD079F13C;	14'h0D02: data <= 32'hD0550244;	14'h0D03: data <= 32'hD030134D;	14'h0D04: data <= 32'hD00B2456;	14'h0D05: data <= 32'hCFE6355E;	14'h0D06: data <= 32'hCFBCA46A;	14'h0D07: data <= 32'hCF90C277;	14'h0D08: data <= 32'hCF64E084;	14'h0D09: data <= 32'hCF38FE90;	14'h0D0A: data <= 32'hCF0D1C9D;	14'h0D0B: data <= 32'hCEE13AAA;	14'h0D0C: data <= 32'hCEB558B7;	14'h0D0D: data <= 32'hCE8976C4;	14'h0D0E: data <= 32'hCE5D94D1;	14'h0D0F: data <= 32'hCE31B2DE;	14'h0D10: data <= 32'hCE05D0EB;	14'h0D11: data <= 32'hCDD9EEF8;	14'h0D12: data <= 32'hCDAE0D05;	14'h0D13: data <= 32'hCD822B12;	14'h0D14: data <= 32'hCD56491E;	14'h0D15: data <= 32'hCD2A672B;	14'h0D16: data <= 32'hCCFE8538;	14'h0D17: data <= 32'hCCD2A345;	14'h0D18: data <= 32'hCCA6C152;	14'h0D19: data <= 32'hCC7ADF5F;	14'h0D1A: data <= 32'hCC4EFD6C;	14'h0D1B: data <= 32'hCC231B79;	14'h0D1C: data <= 32'hCBF73986;	14'h0D1D: data <= 32'hCBCB5793;	14'h0D1E: data <= 32'hCB9F759F;	14'h0D1F: data <= 32'hCB7393AC;	14'h0D20: data <= 32'hCB47B1B9;	14'h0D21: data <= 32'hCB1BCFC6;	14'h0D22: data <= 32'hCAEFEDD3;	14'h0D23: data <= 32'hCAC40BE0;	14'h0D24: data <= 32'hCA95CAF4;	14'h0D25: data <= 32'hCA6363D6;	14'h0D26: data <= 32'hCA30FCB8;	14'h0D27: data <= 32'hC9FE9599;	14'h0D28: data <= 32'hC9CC2E7B;	14'h0D29: data <= 32'hC999C75C;	14'h0D2A: data <= 32'hC967603E;	14'h0D2B: data <= 32'hC934F91F;	14'h0D2C: data <= 32'hC9029201;	14'h0D2D: data <= 32'hC8D02AE2;	14'h0D2E: data <= 32'hC89DC3C4;	14'h0D2F: data <= 32'hC86B5CA5;	14'h0D30: data <= 32'hC838F587;	14'h0D31: data <= 32'hC8068E68;	14'h0D32: data <= 32'hC7D4274A;	14'h0D33: data <= 32'hC7A1C02C;	14'h0D34: data <= 32'hC76F590D;	14'h0D35: data <= 32'hC73CF1EF;	14'h0D36: data <= 32'hC70A8AD0;	14'h0D37: data <= 32'hC6D823B2;	14'h0D38: data <= 32'hC6A5BC93;	14'h0D39: data <= 32'hC6735575;	14'h0D3A: data <= 32'hC640EE56;	14'h0D3B: data <= 32'hC60E8738;	14'h0D3C: data <= 32'hC5DC2019;	14'h0D3D: data <= 32'hC5A9B8FB;	14'h0D3E: data <= 32'hC57751DC;	14'h0D3F: data <= 32'hC544EABE;	14'h0D40: data <= 32'hC51283A0;	14'h0D41: data <= 32'hC4E01C81;	14'h0D42: data <= 32'hC4AD7081;	14'h0D43: data <= 32'hC47698D0;	14'h0D44: data <= 32'hC43FC11E;	14'h0D45: data <= 32'hC408E96D;	14'h0D46: data <= 32'hC3D211BC;	14'h0D47: data <= 32'hC39B3A0B;	14'h0D48: data <= 32'hC364625A;	14'h0D49: data <= 32'hC32D8AA9;	14'h0D4A: data <= 32'hC2F6B2F8;	14'h0D4B: data <= 32'hC2BFDB47;	14'h0D4C: data <= 32'hC2890396;	14'h0D4D: data <= 32'hC2522BE5;	14'h0D4E: data <= 32'hC21B5434;	14'h0D4F: data <= 32'hC1E47C83;	14'h0D50: data <= 32'hC1ADA4D2;	14'h0D51: data <= 32'hC176CD21;	14'h0D52: data <= 32'hC13FF570;	14'h0D53: data <= 32'hC1091DBF;	14'h0D54: data <= 32'hC0D2460E;	14'h0D55: data <= 32'hC09B6E5D;	14'h0D56: data <= 32'hC06496AC;	14'h0D57: data <= 32'hC02DBEFB;	14'h0D58: data <= 32'hBFF6E74A;	14'h0D59: data <= 32'hBFC00F99;	14'h0D5A: data <= 32'hBF8937E8;	14'h0D5B: data <= 32'hBF526036;	14'h0D5C: data <= 32'hBF1B8885;	14'h0D5D: data <= 32'hBEE4B0D4;	14'h0D5E: data <= 32'hBEADD923;	14'h0D5F: data <= 32'hBE770172;	14'h0D60: data <= 32'hBE4029C1;	14'h0D61: data <= 32'hBE08C4A3;	14'h0D62: data <= 32'hBDD13243;	14'h0D63: data <= 32'hBD999FE3;	14'h0D64: data <= 32'hBD620D83;	14'h0D65: data <= 32'hBD2A7B23;	14'h0D66: data <= 32'hBCF2E8C3;	14'h0D67: data <= 32'hBCBB5663;	14'h0D68: data <= 32'hBC83C403;	14'h0D69: data <= 32'hBC4C31A3;	14'h0D6A: data <= 32'hBC149F43;	14'h0D6B: data <= 32'hBBDD0CE3;	14'h0D6C: data <= 32'hBBA57A83;	14'h0D6D: data <= 32'hBB6DE823;	14'h0D6E: data <= 32'hBB3655C3;	14'h0D6F: data <= 32'hBAFEC363;	14'h0D70: data <= 32'hBAC73103;	14'h0D71: data <= 32'hBA8F9EA3;	14'h0D72: data <= 32'hBA580C43;	14'h0D73: data <= 32'hBA2079E3;	14'h0D74: data <= 32'hB9E8E783;	14'h0D75: data <= 32'hB9B15523;	14'h0D76: data <= 32'hB979C2C3;	14'h0D77: data <= 32'hB9423063;	14'h0D78: data <= 32'hB90A9E03;	14'h0D79: data <= 32'hB8D30BA3;	14'h0D7A: data <= 32'hB89B7943;	14'h0D7B: data <= 32'hB863E6E3;	14'h0D7C: data <= 32'hB82C5483;	14'h0D7D: data <= 32'hB7F4C223;	14'h0D7E: data <= 32'hB7BD2FC3;	14'h0D7F: data <= 32'hB7871141;	14'h0D80: data <= 32'hB752B0FE;	14'h0D81: data <= 32'hB71E50BB;	14'h0D82: data <= 32'hB6E9F078;	14'h0D83: data <= 32'hB6B59035;	14'h0D84: data <= 32'hB6812FF2;	14'h0D85: data <= 32'hB64CCFAE;	14'h0D86: data <= 32'hB6186F6B;	14'h0D87: data <= 32'hB5E40F28;	14'h0D88: data <= 32'hB5AFAEE5;	14'h0D89: data <= 32'hB57B4EA2;	14'h0D8A: data <= 32'hB546EE5F;	14'h0D8B: data <= 32'hB5128E1B;	14'h0D8C: data <= 32'hB4DE2DD8;	14'h0D8D: data <= 32'hB4A9CD95;	14'h0D8E: data <= 32'hB4756D52;	14'h0D8F: data <= 32'hB4410D0F;	14'h0D90: data <= 32'hB40CACCC;	14'h0D91: data <= 32'hB3D84C88;	14'h0D92: data <= 32'hB3A3EC45;	14'h0D93: data <= 32'hB36F8C02;	14'h0D94: data <= 32'hB33B2BBF;	14'h0D95: data <= 32'hB306CB7C;	14'h0D96: data <= 32'hB2D26B39;	14'h0D97: data <= 32'hB29E0AF5;	14'h0D98: data <= 32'hB269AAB2;	14'h0D99: data <= 32'hB2354A6F;	14'h0D9A: data <= 32'hB200EA2C;	14'h0D9B: data <= 32'hB1CC89E9;	14'h0D9C: data <= 32'hB19829A6;	14'h0D9D: data <= 32'hB164B5A7;	14'h0D9E: data <= 32'hB1366CBE;	14'h0D9F: data <= 32'hB10823D6;	14'h0DA0: data <= 32'hB0D9DAEE;	14'h0DA1: data <= 32'hB0AB9206;	14'h0DA2: data <= 32'hB07D491E;	14'h0DA3: data <= 32'hB04F0036;	14'h0DA4: data <= 32'hB020B74E;	14'h0DA5: data <= 32'hAFF26E66;	14'h0DA6: data <= 32'hAFC4257E;	14'h0DA7: data <= 32'hAF95DC96;	14'h0DA8: data <= 32'hAF6793AD;	14'h0DA9: data <= 32'hAF394AC5;	14'h0DAA: data <= 32'hAF0B01DD;	14'h0DAB: data <= 32'hAEDCB8F5;	14'h0DAC: data <= 32'hAEAE700D;	14'h0DAD: data <= 32'hAE802725;	14'h0DAE: data <= 32'hAE51DE3D;	14'h0DAF: data <= 32'hAE239555;	14'h0DB0: data <= 32'hADF54C6D;	14'h0DB1: data <= 32'hADC70384;	14'h0DB2: data <= 32'hAD98BA9C;	14'h0DB3: data <= 32'hAD6A71B4;	14'h0DB4: data <= 32'hAD3C28CC;	14'h0DB5: data <= 32'hAD0DDFE4;	14'h0DB6: data <= 32'hACDF96FC;	14'h0DB7: data <= 32'hACB14E14;	14'h0DB8: data <= 32'hAC83052C;	14'h0DB9: data <= 32'hAC54BC44;	14'h0DBA: data <= 32'hAC26735C;	14'h0DBB: data <= 32'hABF82A73;	14'h0DBC: data <= 32'hABD0F5CE;	14'h0DBD: data <= 32'hABAB04C7;	14'h0DBE: data <= 32'hAB8513BF;	14'h0DBF: data <= 32'hAB5F22B8;	14'h0DC0: data <= 32'hAB3931B0;	14'h0DC1: data <= 32'hAB1340A9;	14'h0DC2: data <= 32'hAAED4FA2;	14'h0DC3: data <= 32'hAAC75E9A;	14'h0DC4: data <= 32'hAAA16D93;	14'h0DC5: data <= 32'hAA7B7C8B;	14'h0DC6: data <= 32'hAA558B84;	14'h0DC7: data <= 32'hAA2F9A7D;	14'h0DC8: data <= 32'hAA09A975;	14'h0DC9: data <= 32'hA9E3B86E;	14'h0DCA: data <= 32'hA9BDC767;	14'h0DCB: data <= 32'hA997D65F;	14'h0DCC: data <= 32'hA971E558;	14'h0DCD: data <= 32'hA94BF450;	14'h0DCE: data <= 32'hA9260349;	14'h0DCF: data <= 32'hA9001242;	14'h0DD0: data <= 32'hA8DA213A;	14'h0DD1: data <= 32'hA8B43033;	14'h0DD2: data <= 32'hA88E3F2C;	14'h0DD3: data <= 32'hA8684E24;	14'h0DD4: data <= 32'hA8425D1D;	14'h0DD5: data <= 32'hA81C6C15;	14'h0DD6: data <= 32'hA7F67B0E;	14'h0DD7: data <= 32'hA7D08A07;	14'h0DD8: data <= 32'hA7AA98FF;	14'h0DD9: data <= 32'hA784A7F8;	14'h0DDA: data <= 32'hA7647572;	14'h0DDB: data <= 32'hA7490C58;	14'h0DDC: data <= 32'hA72DA33F;	14'h0DDD: data <= 32'hA7123A25;	14'h0DDE: data <= 32'hA6F6D10B;	14'h0DDF: data <= 32'hA6DB67F2;	14'h0DE0: data <= 32'hA6BFFED8;	14'h0DE1: data <= 32'hA6A495BE;	14'h0DE2: data <= 32'hA6892CA4;	14'h0DE3: data <= 32'hA66DC38B;	14'h0DE4: data <= 32'hA6525A71;	14'h0DE5: data <= 32'hA636F157;	14'h0DE6: data <= 32'hA61B883E;	14'h0DE7: data <= 32'hA6001F24;	14'h0DE8: data <= 32'hA5E4B60A;	14'h0DE9: data <= 32'hA5C94CF1;	14'h0DEA: data <= 32'hA5ADE3D7;	14'h0DEB: data <= 32'hA5927ABD;	14'h0DEC: data <= 32'hA57711A3;	14'h0DED: data <= 32'hA55BA88A;	14'h0DEE: data <= 32'hA5403F70;	14'h0DEF: data <= 32'hA524D656;	14'h0DF0: data <= 32'hA5096D3D;	14'h0DF1: data <= 32'hA4EE0423;	14'h0DF2: data <= 32'hA4D29B09;	14'h0DF3: data <= 32'hA4B731F0;	14'h0DF4: data <= 32'hA49BC8D6;	14'h0DF5: data <= 32'hA4805FBC;	14'h0DF6: data <= 32'hA464F6A2;	14'h0DF7: data <= 32'hA4498D89;	14'h0DF8: data <= 32'hA430EB3A;	14'h0DF9: data <= 32'hA420F628;	14'h0DFA: data <= 32'hA4110115;	14'h0DFB: data <= 32'hA4010C03;	14'h0DFC: data <= 32'hA3F116F0;	14'h0DFD: data <= 32'hA3E121DE;	14'h0DFE: data <= 32'hA3D12CCB;	14'h0DFF: data <= 32'hA3C137B8;	14'h0E00: data <= 32'hA3B142A6;	14'h0E01: data <= 32'hA3A14D93;	14'h0E02: data <= 32'hA3915881;	14'h0E03: data <= 32'hA381636E;	14'h0E04: data <= 32'hA3716E5B;	14'h0E05: data <= 32'hA3617949;	14'h0E06: data <= 32'hA3518436;	14'h0E07: data <= 32'hA3418F24;	14'h0E08: data <= 32'hA3319A11;	14'h0E09: data <= 32'hA321A4FF;	14'h0E0A: data <= 32'hA311AFEC;	14'h0E0B: data <= 32'hA301BAD9;	14'h0E0C: data <= 32'hA2F1C5C7;	14'h0E0D: data <= 32'hA2E1D0B4;	14'h0E0E: data <= 32'hA2D1DBA2;	14'h0E0F: data <= 32'hA2C1E68F;	14'h0E10: data <= 32'hA2B1F17C;	14'h0E11: data <= 32'hA2A1FC6A;	14'h0E12: data <= 32'hA2920757;	14'h0E13: data <= 32'hA2821245;	14'h0E14: data <= 32'hA2721D32;	14'h0E15: data <= 32'hA2622820;	14'h0E16: data <= 32'hA252330D;	14'h0E17: data <= 32'hA24BE49F;	14'h0E18: data <= 32'hA2463597;	14'h0E19: data <= 32'hA240868F;	14'h0E1A: data <= 32'hA23AD786;	14'h0E1B: data <= 32'hA235287E;	14'h0E1C: data <= 32'hA22F7976;	14'h0E1D: data <= 32'hA229CA6D;	14'h0E1E: data <= 32'hA2241B65;	14'h0E1F: data <= 32'hA21E6C5D;	14'h0E20: data <= 32'hA218BD54;	14'h0E21: data <= 32'hA2130E4C;	14'h0E22: data <= 32'hA20D5F44;	14'h0E23: data <= 32'hA207B03B;	14'h0E24: data <= 32'hA2020133;	14'h0E25: data <= 32'hA1FC522B;	14'h0E26: data <= 32'hA1F6A322;	14'h0E27: data <= 32'hA1F0F41A;	14'h0E28: data <= 32'hA1EB4512;	14'h0E29: data <= 32'hA1E59609;	14'h0E2A: data <= 32'hA1DFE701;	14'h0E2B: data <= 32'hA1DA37F9;	14'h0E2C: data <= 32'hA1D488F0;	14'h0E2D: data <= 32'hA1CED9E8;	14'h0E2E: data <= 32'hA1C92AE0;	14'h0E2F: data <= 32'hA1C37BD7;	14'h0E30: data <= 32'hA1BDCCCF;	14'h0E31: data <= 32'hA1B81DC7;	14'h0E32: data <= 32'hA1B26EBE;	14'h0E33: data <= 32'hA1ACBFB6;	14'h0E34: data <= 32'hA1A710AE;	14'h0E35: data <= 32'hA1A6836B;	14'h0E36: data <= 32'hA1A8E4E3;	14'h0E37: data <= 32'hA1AB465A;	14'h0E38: data <= 32'hA1ADA7D1;	14'h0E39: data <= 32'hA1B00949;	14'h0E3A: data <= 32'hA1B26AC0;	14'h0E3B: data <= 32'hA1B4CC38;	14'h0E3C: data <= 32'hA1B72DAF;	14'h0E3D: data <= 32'hA1B98F26;	14'h0E3E: data <= 32'hA1BBF09E;	14'h0E3F: data <= 32'hA1BE5215;	14'h0E40: data <= 32'hA1C0B38D;	14'h0E41: data <= 32'hA1C31504;	14'h0E42: data <= 32'hA1C5767B;	14'h0E43: data <= 32'hA1C7D7F3;	14'h0E44: data <= 32'hA1CA396A;	14'h0E45: data <= 32'hA1CC9AE2;	14'h0E46: data <= 32'hA1CEFC59;	14'h0E47: data <= 32'hA1D15DD0;	14'h0E48: data <= 32'hA1D3BF48;	14'h0E49: data <= 32'hA1D620BF;	14'h0E4A: data <= 32'hA1D88237;	14'h0E4B: data <= 32'hA1DAE3AE;	14'h0E4C: data <= 32'hA1DD4525;	14'h0E4D: data <= 32'hA1DFA69D;	14'h0E4E: data <= 32'hA1E20814;	14'h0E4F: data <= 32'hA1E4698C;	14'h0E50: data <= 32'hA1E6CB03;	14'h0E51: data <= 32'hA1E92C7A;	14'h0E52: data <= 32'hA1EB8DF2;	14'h0E53: data <= 32'hA1F00EFD;	14'h0E54: data <= 32'hA1F8CF31;	14'h0E55: data <= 32'hA2018F64;	14'h0E56: data <= 32'hA20A4F98;	14'h0E57: data <= 32'hA2130FCB;	14'h0E58: data <= 32'hA21BCFFF;	14'h0E59: data <= 32'hA2249032;	14'h0E5A: data <= 32'hA22D5066;	14'h0E5B: data <= 32'hA2361099;	14'h0E5C: data <= 32'hA23ED0CD;	14'h0E5D: data <= 32'hA2479100;	14'h0E5E: data <= 32'hA2505134;	14'h0E5F: data <= 32'hA2591167;	14'h0E60: data <= 32'hA261D19B;	14'h0E61: data <= 32'hA26A91CE;	14'h0E62: data <= 32'hA2735202;	14'h0E63: data <= 32'hA27C1235;	14'h0E64: data <= 32'hA284D269;	14'h0E65: data <= 32'hA28D929C;	14'h0E66: data <= 32'hA29652D0;	14'h0E67: data <= 32'hA29F1303;	14'h0E68: data <= 32'hA2A7D337;	14'h0E69: data <= 32'hA2B0936A;	14'h0E6A: data <= 32'hA2B9539E;	14'h0E6B: data <= 32'hA2C213D1;	14'h0E6C: data <= 32'hA2CAD405;	14'h0E6D: data <= 32'hA2D39438;	14'h0E6E: data <= 32'hA2DC546C;	14'h0E6F: data <= 32'hA2E5149F;	14'h0E70: data <= 32'hA2EDD4D3;	14'h0E71: data <= 32'hA2F6B7F7;	14'h0E72: data <= 32'hA303F936;	14'h0E73: data <= 32'hA3113A75;	14'h0E74: data <= 32'hA31E7BB4;	14'h0E75: data <= 32'hA32BBCF3;	14'h0E76: data <= 32'hA338FE31;	14'h0E77: data <= 32'hA3463F70;	14'h0E78: data <= 32'hA35380AF;	14'h0E79: data <= 32'hA360C1EE;	14'h0E7A: data <= 32'hA36E032D;	14'h0E7B: data <= 32'hA37B446C;	14'h0E7C: data <= 32'hA38885AB;	14'h0E7D: data <= 32'hA395C6EA;	14'h0E7E: data <= 32'hA3A30829;	14'h0E7F: data <= 32'hA3B04968;	14'h0E80: data <= 32'hA3BD8AA7;	14'h0E81: data <= 32'hA3CACBE5;	14'h0E82: data <= 32'hA3D80D24;	14'h0E83: data <= 32'hA3E54E63;	14'h0E84: data <= 32'hA3F28FA2;	14'h0E85: data <= 32'hA3FFD0E1;	14'h0E86: data <= 32'hA40D1220;	14'h0E87: data <= 32'hA41A535F;	14'h0E88: data <= 32'hA427949E;	14'h0E89: data <= 32'hA434D5DD;	14'h0E8A: data <= 32'hA442171C;	14'h0E8B: data <= 32'hA44F585B;	14'h0E8C: data <= 32'hA45C999A;	14'h0E8D: data <= 32'hA469DAD8;	14'h0E8E: data <= 32'hA4771C17;	14'h0E8F: data <= 32'hA4845D56;	14'h0E90: data <= 32'hA49315F2;	14'h0E91: data <= 32'hA4A25B51;	14'h0E92: data <= 32'hA4B1A0B0;	14'h0E93: data <= 32'hA4C0E60F;	14'h0E94: data <= 32'hA4D02B6E;	14'h0E95: data <= 32'hA4DF70CC;	14'h0E96: data <= 32'hA4EEB62B;	14'h0E97: data <= 32'hA4FDFB8A;	14'h0E98: data <= 32'hA50D40E9;	14'h0E99: data <= 32'hA51C8648;	14'h0E9A: data <= 32'hA52BCBA7;	14'h0E9B: data <= 32'hA53B1106;	14'h0E9C: data <= 32'hA54A5664;	14'h0E9D: data <= 32'hA5599BC3;	14'h0E9E: data <= 32'hA568E122;	14'h0E9F: data <= 32'hA5782681;	14'h0EA0: data <= 32'hA5876BE0;	14'h0EA1: data <= 32'hA596B13F;	14'h0EA2: data <= 32'hA5A5F69E;	14'h0EA3: data <= 32'hA5B53BFC;	14'h0EA4: data <= 32'hA5C4815B;	14'h0EA5: data <= 32'hA5D3C6BA;	14'h0EA6: data <= 32'hA5E30C19;	14'h0EA7: data <= 32'hA5F25178;	14'h0EA8: data <= 32'hA60196D7;	14'h0EA9: data <= 32'hA610DC36;	14'h0EAA: data <= 32'hA6202194;	14'h0EAB: data <= 32'hA62F66F3;	14'h0EAC: data <= 32'hA63EAC52;	14'h0EAD: data <= 32'hA64DF1B1;	14'h0EAE: data <= 32'hA65D1FC5;	14'h0EAF: data <= 32'hA66C2E3B;	14'h0EB0: data <= 32'hA67B3CB2;	14'h0EB1: data <= 32'hA68A4B29;	14'h0EB2: data <= 32'hA699599F;	14'h0EB3: data <= 32'hA6A86816;	14'h0EB4: data <= 32'hA6B7768D;	14'h0EB5: data <= 32'hA6C68503;	14'h0EB6: data <= 32'hA6D5937A;	14'h0EB7: data <= 32'hA6E4A1F1;	14'h0EB8: data <= 32'hA6F3B067;	14'h0EB9: data <= 32'hA702BEDE;	14'h0EBA: data <= 32'hA711CD55;	14'h0EBB: data <= 32'hA720DBCB;	14'h0EBC: data <= 32'hA72FEA42;	14'h0EBD: data <= 32'hA73EF8B9;	14'h0EBE: data <= 32'hA74E072F;	14'h0EBF: data <= 32'hA75D15A6;	14'h0EC0: data <= 32'hA76C241D;	14'h0EC1: data <= 32'hA77B3293;	14'h0EC2: data <= 32'hA78A410A;	14'h0EC3: data <= 32'hA7994F81;	14'h0EC4: data <= 32'hA7A85DF7;	14'h0EC5: data <= 32'hA7B76C6E;	14'h0EC6: data <= 32'hA7C67AE5;	14'h0EC7: data <= 32'hA7D5895B;	14'h0EC8: data <= 32'hA7E497D2;	14'h0EC9: data <= 32'hA7F3A649;	14'h0ECA: data <= 32'hA802B4BF;	14'h0ECB: data <= 32'hA811C336;	14'h0ECC: data <= 32'hA820A9BE;	14'h0ECD: data <= 32'hA82E6EC4;	14'h0ECE: data <= 32'hA83C33C9;	14'h0ECF: data <= 32'hA849F8CF;	14'h0ED0: data <= 32'hA857BDD5;	14'h0ED1: data <= 32'hA86582DB;	14'h0ED2: data <= 32'hA87347E0;	14'h0ED3: data <= 32'hA8810CE6;	14'h0ED4: data <= 32'hA88ED1EC;	14'h0ED5: data <= 32'hA89C96F2;	14'h0ED6: data <= 32'hA8AA5BF7;	14'h0ED7: data <= 32'hA8B820FD;	14'h0ED8: data <= 32'hA8C5E603;	14'h0ED9: data <= 32'hA8D3AB08;	14'h0EDA: data <= 32'hA8E1700E;	14'h0EDB: data <= 32'hA8EF3514;	14'h0EDC: data <= 32'hA8FCFA1A;	14'h0EDD: data <= 32'hA90ABF1F;	14'h0EDE: data <= 32'hA9188425;	14'h0EDF: data <= 32'hA926492B;	14'h0EE0: data <= 32'hA9340E30;	14'h0EE1: data <= 32'hA941D336;	14'h0EE2: data <= 32'hA94F983C;	14'h0EE3: data <= 32'hA95D5D42;	14'h0EE4: data <= 32'hA96B2247;	14'h0EE5: data <= 32'hA978E74D;	14'h0EE6: data <= 32'hA986AC53;	14'h0EE7: data <= 32'hA9947159;	14'h0EE8: data <= 32'hA9A2365E;	14'h0EE9: data <= 32'hA9AFFB64;	14'h0EEA: data <= 32'hA9BDC06A;	14'h0EEB: data <= 32'hA9C9F59D;	14'h0EEC: data <= 32'hA9D5D1F7;	14'h0EED: data <= 32'hA9E1AE51;	14'h0EEE: data <= 32'hA9ED8AAB;	14'h0EEF: data <= 32'hA9F96704;	14'h0EF0: data <= 32'hAA05435E;	14'h0EF1: data <= 32'hAA111FB8;	14'h0EF2: data <= 32'hAA1CFC12;	14'h0EF3: data <= 32'hAA28D86C;	14'h0EF4: data <= 32'hAA34B4C6;	14'h0EF5: data <= 32'hAA409120;	14'h0EF6: data <= 32'hAA4C6D79;	14'h0EF7: data <= 32'hAA5849D3;	14'h0EF8: data <= 32'hAA64262D;	14'h0EF9: data <= 32'hAA700287;	14'h0EFA: data <= 32'hAA7BDEE1;	14'h0EFB: data <= 32'hAA87BB3B;	14'h0EFC: data <= 32'hAA939795;	14'h0EFD: data <= 32'hAA9F73EE;	14'h0EFE: data <= 32'hAAAB5048;	14'h0EFF: data <= 32'hAAB72CA2;	14'h0F00: data <= 32'hAAC308FC;	14'h0F01: data <= 32'hAACEE556;	14'h0F02: data <= 32'hAADAC1B0;	14'h0F03: data <= 32'hAAE69E0A;	14'h0F04: data <= 32'hAAF27A63;	14'h0F05: data <= 32'hAAFE56BD;	14'h0F06: data <= 32'hAB0A3317;	14'h0F07: data <= 32'hAB160F71;	14'h0F08: data <= 32'hAB21EBCB;	14'h0F09: data <= 32'hAB2C74B8;	14'h0F0A: data <= 32'hAB35BE30;	14'h0F0B: data <= 32'hAB3F07A8;	14'h0F0C: data <= 32'hAB485120;	14'h0F0D: data <= 32'hAB519A98;	14'h0F0E: data <= 32'hAB5AE40F;	14'h0F0F: data <= 32'hAB642D87;	14'h0F10: data <= 32'hAB6D76FF;	14'h0F11: data <= 32'hAB76C077;	14'h0F12: data <= 32'hAB8009EF;	14'h0F13: data <= 32'hAB895367;	14'h0F14: data <= 32'hAB929CDF;	14'h0F15: data <= 32'hAB9BE657;	14'h0F16: data <= 32'hABA52FCE;	14'h0F17: data <= 32'hABAE7946;	14'h0F18: data <= 32'hABB7C2BE;	14'h0F19: data <= 32'hABC10C36;	14'h0F1A: data <= 32'hABCA55AE;	14'h0F1B: data <= 32'hABD39F26;	14'h0F1C: data <= 32'hABDCE89E;	14'h0F1D: data <= 32'hABE63216;	14'h0F1E: data <= 32'hABEF7B8D;	14'h0F1F: data <= 32'hABF8C505;	14'h0F20: data <= 32'hAC020E7D;	14'h0F21: data <= 32'hAC0B57F5;	14'h0F22: data <= 32'hAC14A16D;	14'h0F23: data <= 32'hAC1DEAE5;	14'h0F24: data <= 32'hAC27345D;	14'h0F25: data <= 32'hAC307DD4;	14'h0F26: data <= 32'hAC39C74C;	14'h0F27: data <= 32'hAC42725E;	14'h0F28: data <= 32'hAC48D11A;	14'h0F29: data <= 32'hAC4F2FD6;	14'h0F2A: data <= 32'hAC558E92;	14'h0F2B: data <= 32'hAC5BED4F;	14'h0F2C: data <= 32'hAC624C0B;	14'h0F2D: data <= 32'hAC68AAC7;	14'h0F2E: data <= 32'hAC6F0983;	14'h0F2F: data <= 32'hAC75683F;	14'h0F30: data <= 32'hAC7BC6FB;	14'h0F31: data <= 32'hAC8225B7;	14'h0F32: data <= 32'hAC888473;	14'h0F33: data <= 32'hAC8EE32F;	14'h0F34: data <= 32'hAC9541EB;	14'h0F35: data <= 32'hAC9BA0A7;	14'h0F36: data <= 32'hACA1FF63;	14'h0F37: data <= 32'hACA85E1F;	14'h0F38: data <= 32'hACAEBCDB;	14'h0F39: data <= 32'hACB51B97;	14'h0F3A: data <= 32'hACBB7A53;	14'h0F3B: data <= 32'hACC1D90F;	14'h0F3C: data <= 32'hACC837CB;	14'h0F3D: data <= 32'hACCE9687;	14'h0F3E: data <= 32'hACD4F544;	14'h0F3F: data <= 32'hACDB5400;	14'h0F40: data <= 32'hACE1B2BC;	14'h0F41: data <= 32'hACE81178;	14'h0F42: data <= 32'hACEE7034;	14'h0F43: data <= 32'hACF4CEF0;	14'h0F44: data <= 32'hACFB2DAC;	14'h0F45: data <= 32'hAD018C68;	14'h0F46: data <= 32'hAD05EE01;	14'h0F47: data <= 32'hAD0A1CB0;	14'h0F48: data <= 32'hAD0E4B5F;	14'h0F49: data <= 32'hAD127A0F;	14'h0F4A: data <= 32'hAD16A8BE;	14'h0F4B: data <= 32'hAD1AD76D;	14'h0F4C: data <= 32'hAD1F061C;	14'h0F4D: data <= 32'hAD2334CB;	14'h0F4E: data <= 32'hAD27637B;	14'h0F4F: data <= 32'hAD2B922A;	14'h0F50: data <= 32'hAD2FC0D9;	14'h0F51: data <= 32'hAD33EF88;	14'h0F52: data <= 32'hAD381E37;	14'h0F53: data <= 32'hAD3C4CE6;	14'h0F54: data <= 32'hAD407B96;	14'h0F55: data <= 32'hAD44AA45;	14'h0F56: data <= 32'hAD48D8F4;	14'h0F57: data <= 32'hAD4D07A3;	14'h0F58: data <= 32'hAD513652;	14'h0F59: data <= 32'hAD556502;	14'h0F5A: data <= 32'hAD5993B1;	14'h0F5B: data <= 32'hAD5DC260;	14'h0F5C: data <= 32'hAD61F10F;	14'h0F5D: data <= 32'hAD661FBE;	14'h0F5E: data <= 32'hAD6A4E6E;	14'h0F5F: data <= 32'hAD6E7D1D;	14'h0F60: data <= 32'hAD72ABCC;	14'h0F61: data <= 32'hAD76DA7B;	14'h0F62: data <= 32'hAD7B092A;	14'h0F63: data <= 32'hAD7F37DA;	14'h0F64: data <= 32'hAD830CB0;	14'h0F65: data <= 32'hAD86A71F;	14'h0F66: data <= 32'hAD8A418F;	14'h0F67: data <= 32'hAD8DDBFE;	14'h0F68: data <= 32'hAD91766E;	14'h0F69: data <= 32'hAD9510DE;	14'h0F6A: data <= 32'hAD98AB4D;	14'h0F6B: data <= 32'hAD9C45BD;	14'h0F6C: data <= 32'hAD9FE02C;	14'h0F6D: data <= 32'hADA37A9C;	14'h0F6E: data <= 32'hADA7150B;	14'h0F6F: data <= 32'hADAAAF7B;	14'h0F70: data <= 32'hADAE49EA;	14'h0F71: data <= 32'hADB1E45A;	14'h0F72: data <= 32'hADB57EC9;	14'h0F73: data <= 32'hADB91939;	14'h0F74: data <= 32'hADBCB3A9;	14'h0F75: data <= 32'hADC04E18;	14'h0F76: data <= 32'hADC3E888;	14'h0F77: data <= 32'hADC782F7;	14'h0F78: data <= 32'hADCB1D67;	14'h0F79: data <= 32'hADCEB7D6;	14'h0F7A: data <= 32'hADD25246;	14'h0F7B: data <= 32'hADD5ECB5;	14'h0F7C: data <= 32'hADD98725;	14'h0F7D: data <= 32'hADDD2194;	14'h0F7E: data <= 32'hADE0BC04;	14'h0F7F: data <= 32'hADE45674;	14'h0F80: data <= 32'hADE7F0E3;	14'h0F81: data <= 32'hADEB8B53;	14'h0F82: data <= 32'hADEF7C47;	14'h0F83: data <= 32'hADF4343B;	14'h0F84: data <= 32'hADF8EC2E;	14'h0F85: data <= 32'hADFDA422;	14'h0F86: data <= 32'hAE025C16;	14'h0F87: data <= 32'hAE071409;	14'h0F88: data <= 32'hAE0BCBFD;	14'h0F89: data <= 32'hAE1083F1;	14'h0F8A: data <= 32'hAE153BE4;	14'h0F8B: data <= 32'hAE19F3D8;	14'h0F8C: data <= 32'hAE1EABCB;	14'h0F8D: data <= 32'hAE2363BF;	14'h0F8E: data <= 32'hAE281BB3;	14'h0F8F: data <= 32'hAE2CD3A6;	14'h0F90: data <= 32'hAE318B9A;	14'h0F91: data <= 32'hAE36438D;	14'h0F92: data <= 32'hAE3AFB81;	14'h0F93: data <= 32'hAE3FB375;	14'h0F94: data <= 32'hAE446B68;	14'h0F95: data <= 32'hAE49235C;	14'h0F96: data <= 32'hAE4DDB4F;	14'h0F97: data <= 32'hAE529343;	14'h0F98: data <= 32'hAE574B37;	14'h0F99: data <= 32'hAE5C032A;	14'h0F9A: data <= 32'hAE60BB1E;	14'h0F9B: data <= 32'hAE657311;	14'h0F9C: data <= 32'hAE6A2B05;	14'h0F9D: data <= 32'hAE6EE2F9;	14'h0F9E: data <= 32'hAE739AEC;	14'h0F9F: data <= 32'hAE7852E0;	14'h0FA0: data <= 32'hAE7D0AD3;	14'h0FA1: data <= 32'hAE84711D;	14'h0FA2: data <= 32'hAE8BD767;	14'h0FA3: data <= 32'hAE933DB0;	14'h0FA4: data <= 32'hAE9AA3FA;	14'h0FA5: data <= 32'hAEA20A44;	14'h0FA6: data <= 32'hAEA9708D;	14'h0FA7: data <= 32'hAEB0D6D7;	14'h0FA8: data <= 32'hAEB83D21;	14'h0FA9: data <= 32'hAEBFA36A;	14'h0FAA: data <= 32'hAEC709B4;	14'h0FAB: data <= 32'hAECE6FFE;	14'h0FAC: data <= 32'hAED5D647;	14'h0FAD: data <= 32'hAEDD3C91;	14'h0FAE: data <= 32'hAEE4A2DA;	14'h0FAF: data <= 32'hAEEC0924;	14'h0FB0: data <= 32'hAEF36F6E;	14'h0FB1: data <= 32'hAEFAD5B7;	14'h0FB2: data <= 32'hAF023C01;	14'h0FB3: data <= 32'hAF09A24B;	14'h0FB4: data <= 32'hAF110894;	14'h0FB5: data <= 32'hAF186EDE;	14'h0FB6: data <= 32'hAF1FD528;	14'h0FB7: data <= 32'hAF273B71;	14'h0FB8: data <= 32'hAF2EA1BB;	14'h0FB9: data <= 32'hAF360804;	14'h0FBA: data <= 32'hAF3D6E4E;	14'h0FBB: data <= 32'hAF44D498;	14'h0FBC: data <= 32'hAF4C3AE1;	14'h0FBD: data <= 32'hAF53A12B;	14'h0FBE: data <= 32'hAF5B0775;	14'h0FBF: data <= 32'hAF6531B6;	14'h0FC0: data <= 32'hAF708FC6;	14'h0FC1: data <= 32'hAF7BEDD7;	14'h0FC2: data <= 32'hAF874BE8;	14'h0FC3: data <= 32'hAF92A9F8;	14'h0FC4: data <= 32'hAF9E0809;	14'h0FC5: data <= 32'hAFA9661A;	14'h0FC6: data <= 32'hAFB4C42A;	14'h0FC7: data <= 32'hAFC0223B;	14'h0FC8: data <= 32'hAFCB804C;	14'h0FC9: data <= 32'hAFD6DE5D;	14'h0FCA: data <= 32'hAFE23C6D;	14'h0FCB: data <= 32'hAFED9A7E;	14'h0FCC: data <= 32'hAFF8F88F;	14'h0FCD: data <= 32'hB004569F;	14'h0FCE: data <= 32'hB00FB4B0;	14'h0FCF: data <= 32'hB01B12C1;	14'h0FD0: data <= 32'hB02670D1;	14'h0FD1: data <= 32'hB031CEE2;	14'h0FD2: data <= 32'hB03D2CF3;	14'h0FD3: data <= 32'hB0488B03;	14'h0FD4: data <= 32'hB053E914;	14'h0FD5: data <= 32'hB05F4725;	14'h0FD6: data <= 32'hB06AA535;	14'h0FD7: data <= 32'hB0760346;	14'h0FD8: data <= 32'hB0816157;	14'h0FD9: data <= 32'hB08CBF67;	14'h0FDA: data <= 32'hB0981D78;	14'h0FDB: data <= 32'hB0A37B89;	14'h0FDC: data <= 32'hB0AED999;	14'h0FDD: data <= 32'hB0BC22AA;	14'h0FDE: data <= 32'hB0CC5F1E;	14'h0FDF: data <= 32'hB0DC9B92;	14'h0FE0: data <= 32'hB0ECD805;	14'h0FE1: data <= 32'hB0FD1479;	14'h0FE2: data <= 32'hB10D50EC;	14'h0FE3: data <= 32'hB11D8D60;	14'h0FE4: data <= 32'hB12DC9D4;	14'h0FE5: data <= 32'hB13E0647;	14'h0FE6: data <= 32'hB14E42BB;	14'h0FE7: data <= 32'hB15E7F2E;	14'h0FE8: data <= 32'hB16EBBA2;	14'h0FE9: data <= 32'hB17EF816;	14'h0FEA: data <= 32'hB18F3489;	14'h0FEB: data <= 32'hB19F70FD;	14'h0FEC: data <= 32'hB1AFAD70;	14'h0FED: data <= 32'hB1BFE9E4;	14'h0FEE: data <= 32'hB1D02658;	14'h0FEF: data <= 32'hB1E062CB;	14'h0FF0: data <= 32'hB1F09F3F;	14'h0FF1: data <= 32'hB200DBB2;	14'h0FF2: data <= 32'hB2111826;	14'h0FF3: data <= 32'hB221549A;	14'h0FF4: data <= 32'hB231910D;	14'h0FF5: data <= 32'hB241CD81;	14'h0FF6: data <= 32'hB25209F4;	14'h0FF7: data <= 32'hB2624668;	14'h0FF8: data <= 32'hB27282DC;	14'h0FF9: data <= 32'hB282BF4F;	14'h0FFA: data <= 32'hB292FBC3;	14'h0FFB: data <= 32'hB2A3A607;	14'h0FFC: data <= 32'hB2B89A6E;	14'h0FFD: data <= 32'hB2CD8ED5;	14'h0FFE: data <= 32'hB2E2833C;	14'h0FFF: data <= 32'hB2F777A4;	14'h1000: data <= 32'hB30C6C0B;	14'h1001: data <= 32'hB3216072;	14'h1002: data <= 32'hB33654D9;	14'h1003: data <= 32'hB34B4940;	14'h1004: data <= 32'hB3603DA7;	14'h1005: data <= 32'hB375320F;	14'h1006: data <= 32'hB38A2676;	14'h1007: data <= 32'hB39F1ADD;	14'h1008: data <= 32'hB3B40F44;	14'h1009: data <= 32'hB3C903AB;	14'h100A: data <= 32'hB3DDF812;	14'h100B: data <= 32'hB3F2EC7A;	14'h100C: data <= 32'hB407E0E1;	14'h100D: data <= 32'hB41CD548;	14'h100E: data <= 32'hB431C9AF;	14'h100F: data <= 32'hB446BE16;	14'h1010: data <= 32'hB45BB27E;	14'h1011: data <= 32'hB470A6E5;	14'h1012: data <= 32'hB4859B4C;	14'h1013: data <= 32'hB49A8FB3;	14'h1014: data <= 32'hB4AF841A;	14'h1015: data <= 32'hB4C47881;	14'h1016: data <= 32'hB4D96CE9;	14'h1017: data <= 32'hB4EE6150;	14'h1018: data <= 32'hB50355B7;	14'h1019: data <= 32'hB5184A1E;	14'h101A: data <= 32'hB53051DA;	14'h101B: data <= 32'hB5492D90;	14'h101C: data <= 32'hB5620945;	14'h101D: data <= 32'hB57AE4FA;	14'h101E: data <= 32'hB593C0B0;	14'h101F: data <= 32'hB5AC9C65;	14'h1020: data <= 32'hB5C5781B;	14'h1021: data <= 32'hB5DE53D0;	14'h1022: data <= 32'hB5F72F85;	14'h1023: data <= 32'hB6100B3B;	14'h1024: data <= 32'hB628E6F0;	14'h1025: data <= 32'hB641C2A5;	14'h1026: data <= 32'hB65A9E5B;	14'h1027: data <= 32'hB6737A10;	14'h1028: data <= 32'hB68C55C6;	14'h1029: data <= 32'hB6A5317B;	14'h102A: data <= 32'hB6BE0D30;	14'h102B: data <= 32'hB6D6E8E6;	14'h102C: data <= 32'hB6EFC49B;	14'h102D: data <= 32'hB708A051;	14'h102E: data <= 32'hB7217C06;	14'h102F: data <= 32'hB73A57BB;	14'h1030: data <= 32'hB7533371;	14'h1031: data <= 32'hB76C0F26;	14'h1032: data <= 32'hB784EADB;	14'h1033: data <= 32'hB79DC691;	14'h1034: data <= 32'hB7B6A246;	14'h1035: data <= 32'hB7CF7DFC;	14'h1036: data <= 32'hB7E859B1;	14'h1037: data <= 32'hB8013566;	14'h1038: data <= 32'hB81BA06E;	14'h1039: data <= 32'hB837B3BE;	14'h103A: data <= 32'hB853C70E;	14'h103B: data <= 32'hB86FDA5E;	14'h103C: data <= 32'hB88BEDAE;	14'h103D: data <= 32'hB8A800FD;	14'h103E: data <= 32'hB8C4144D;	14'h103F: data <= 32'hB8E0279D;	14'h1040: data <= 32'hB8FC3AED;	14'h1041: data <= 32'hB9184E3C;	14'h1042: data <= 32'hB934618C;	14'h1043: data <= 32'hB95074DC;	14'h1044: data <= 32'hB96C882C;	14'h1045: data <= 32'hB9889B7C;	14'h1046: data <= 32'hB9A4AECB;	14'h1047: data <= 32'hB9C0C21B;	14'h1048: data <= 32'hB9DCD56B;	14'h1049: data <= 32'hB9F8E8BB;	14'h104A: data <= 32'hBA14FC0B;	14'h104B: data <= 32'hBA310F5A;	14'h104C: data <= 32'hBA4D22AA;	14'h104D: data <= 32'hBA6935FA;	14'h104E: data <= 32'hBA85494A;	14'h104F: data <= 32'hBAA15C9A;	14'h1050: data <= 32'hBABD6FE9;	14'h1051: data <= 32'hBAD98339;	14'h1052: data <= 32'hBAF59689;	14'h1053: data <= 32'hBB11A9D9;	14'h1054: data <= 32'hBB2DBD29;	14'h1055: data <= 32'hBB49D078;	14'h1056: data <= 32'hBB666291;	14'h1057: data <= 32'hBB852F32;	14'h1058: data <= 32'hBBA3FBD3;	14'h1059: data <= 32'hBBC2C875;	14'h105A: data <= 32'hBBE19516;	14'h105B: data <= 32'hBC0061B7;	14'h105C: data <= 32'hBC1F2E58;	14'h105D: data <= 32'hBC3DFAF9;	14'h105E: data <= 32'hBC5CC79A;	14'h105F: data <= 32'hBC7B943B;	14'h1060: data <= 32'hBC9A60DC;	14'h1061: data <= 32'hBCB92D7E;	14'h1062: data <= 32'hBCD7FA1F;	14'h1063: data <= 32'hBCF6C6C0;	14'h1064: data <= 32'hBD159361;	14'h1065: data <= 32'hBD346002;	14'h1066: data <= 32'hBD532CA3;	14'h1067: data <= 32'hBD71F944;	14'h1068: data <= 32'hBD90C5E5;	14'h1069: data <= 32'hBDAF9287;	14'h106A: data <= 32'hBDCE5F28;	14'h106B: data <= 32'hBDED2BC9;	14'h106C: data <= 32'hBE0BF86A;	14'h106D: data <= 32'hBE2AC50B;	14'h106E: data <= 32'hBE4991AC;	14'h106F: data <= 32'hBE685E4D;	14'h1070: data <= 32'hBE872AEF;	14'h1071: data <= 32'hBEA5F790;	14'h1072: data <= 32'hBEC4C431;	14'h1073: data <= 32'hBEE390D2;	14'h1074: data <= 32'hBF025D73;	14'h1075: data <= 32'hBF22AC17;	14'h1076: data <= 32'hBF432FFA;	14'h1077: data <= 32'hBF63B3DC;	14'h1078: data <= 32'hBF8437BE;	14'h1079: data <= 32'hBFA4BBA1;	14'h107A: data <= 32'hBFC53F83;	14'h107B: data <= 32'hBFE5C366;	14'h107C: data <= 32'hC0064748;	14'h107D: data <= 32'hC026CB2B;	14'h107E: data <= 32'hC0474F0D;	14'h107F: data <= 32'hC067D2EF;	14'h1080: data <= 32'hC08856D2;	14'h1081: data <= 32'hC0A8DAB4;	14'h1082: data <= 32'hC0C95E97;	14'h1083: data <= 32'hC0E9E279;	14'h1084: data <= 32'hC10A665B;	14'h1085: data <= 32'hC12AEA3E;	14'h1086: data <= 32'hC14B6E20;	14'h1087: data <= 32'hC16BF203;	14'h1088: data <= 32'hC18C75E5;	14'h1089: data <= 32'hC1ACF9C7;	14'h108A: data <= 32'hC1CD7DAA;	14'h108B: data <= 32'hC1EE018C;	14'h108C: data <= 32'hC20E856F;	14'h108D: data <= 32'hC22F0951;	14'h108E: data <= 32'hC24F8D34;	14'h108F: data <= 32'hC2701116;	14'h1090: data <= 32'hC29094F8;	14'h1091: data <= 32'hC2B118DB;	14'h1092: data <= 32'hC2D19CBD;	14'h1093: data <= 32'hC2F2500B;	14'h1094: data <= 32'hC313264A;	14'h1095: data <= 32'hC333FC88;	14'h1096: data <= 32'hC354D2C7;	14'h1097: data <= 32'hC375A906;	14'h1098: data <= 32'hC3967F44;	14'h1099: data <= 32'hC3B75583;	14'h109A: data <= 32'hC3D82BC1;	14'h109B: data <= 32'hC3F90200;	14'h109C: data <= 32'hC419D83F;	14'h109D: data <= 32'hC43AAE7D;	14'h109E: data <= 32'hC45B84BC;	14'h109F: data <= 32'hC47C5AFB;	14'h10A0: data <= 32'hC49D3139;	14'h10A1: data <= 32'hC4BE0778;	14'h10A2: data <= 32'hC4DEDDB7;	14'h10A3: data <= 32'hC4FFB3F5;	14'h10A4: data <= 32'hC5208A34;	14'h10A5: data <= 32'hC5416073;	14'h10A6: data <= 32'hC56236B1;	14'h10A7: data <= 32'hC5830CF0;	14'h10A8: data <= 32'hC5A3E32E;	14'h10A9: data <= 32'hC5C4B96D;	14'h10AA: data <= 32'hC5E58FAC;	14'h10AB: data <= 32'hC60665EA;	14'h10AC: data <= 32'hC6273C29;	14'h10AD: data <= 32'hC6481268;	14'h10AE: data <= 32'hC668E8A6;	14'h10AF: data <= 32'hC689BEE5;	14'h10B0: data <= 32'hC6AA9524;	14'h10B1: data <= 32'hC6CB2C7E;	14'h10B2: data <= 32'hC6EB1C20;	14'h10B3: data <= 32'hC70B0BC3;	14'h10B4: data <= 32'hC72AFB66;	14'h10B5: data <= 32'hC74AEB09;	14'h10B6: data <= 32'hC76ADAAB;	14'h10B7: data <= 32'hC78ACA4E;	14'h10B8: data <= 32'hC7AAB9F1;	14'h10B9: data <= 32'hC7CAA994;	14'h10BA: data <= 32'hC7EA9936;	14'h10BB: data <= 32'hC80A88D9;	14'h10BC: data <= 32'hC82A787C;	14'h10BD: data <= 32'hC84A681F;	14'h10BE: data <= 32'hC86A57C1;	14'h10BF: data <= 32'hC88A4764;	14'h10C0: data <= 32'hC8AA3707;	14'h10C1: data <= 32'hC8CA26AA;	14'h10C2: data <= 32'hC8EA164C;	14'h10C3: data <= 32'hC90A05EF;	14'h10C4: data <= 32'hC929F592;	14'h10C5: data <= 32'hC949E535;	14'h10C6: data <= 32'hC969D4D8;	14'h10C7: data <= 32'hC989C47A;	14'h10C8: data <= 32'hC9A9B41D;	14'h10C9: data <= 32'hC9C9A3C0;	14'h10CA: data <= 32'hC9E99363;	14'h10CB: data <= 32'hCA098305;	14'h10CC: data <= 32'hCA2972A8;	14'h10CD: data <= 32'hCA49624B;	14'h10CE: data <= 32'hCA6951EE;	14'h10CF: data <= 32'hCA894190;	14'h10D0: data <= 32'hCAA7F711;	14'h10D1: data <= 32'hCAC6A2C0;	14'h10D2: data <= 32'hCAE54E70;	14'h10D3: data <= 32'hCB03FA1F;	14'h10D4: data <= 32'hCB22A5CF;	14'h10D5: data <= 32'hCB41517E;	14'h10D6: data <= 32'hCB5FFD2D;	14'h10D7: data <= 32'hCB7EA8DD;	14'h10D8: data <= 32'hCB9D548C;	14'h10D9: data <= 32'hCBBC003C;	14'h10DA: data <= 32'hCBDAABEB;	14'h10DB: data <= 32'hCBF9579A;	14'h10DC: data <= 32'hCC18034A;	14'h10DD: data <= 32'hCC36AEF9;	14'h10DE: data <= 32'hCC555AA9;	14'h10DF: data <= 32'hCC740658;	14'h10E0: data <= 32'hCC92B208;	14'h10E1: data <= 32'hCCB15DB7;	14'h10E2: data <= 32'hCCD00966;	14'h10E3: data <= 32'hCCEEB516;	14'h10E4: data <= 32'hCD0D60C5;	14'h10E5: data <= 32'hCD2C0C75;	14'h10E6: data <= 32'hCD4AB824;	14'h10E7: data <= 32'hCD6963D4;	14'h10E8: data <= 32'hCD880F83;	14'h10E9: data <= 32'hCDA6BB32;	14'h10EA: data <= 32'hCDC566E2;	14'h10EB: data <= 32'hCDE41291;	14'h10EC: data <= 32'hCE02BE41;	14'h10ED: data <= 32'hCE2169F0;	14'h10EE: data <= 32'hCE3F4C4C;	14'h10EF: data <= 32'hCE5CC9FF;	14'h10F0: data <= 32'hCE7A47B1;	14'h10F1: data <= 32'hCE97C564;	14'h10F2: data <= 32'hCEB54316;	14'h10F3: data <= 32'hCED2C0C9;	14'h10F4: data <= 32'hCEF03E7B;	14'h10F5: data <= 32'hCF0DBC2E;	14'h10F6: data <= 32'hCF2B39E0;	14'h10F7: data <= 32'hCF48B793;	14'h10F8: data <= 32'hCF663545;	14'h10F9: data <= 32'hCF83B2F8;	14'h10FA: data <= 32'hCFA130AA;	14'h10FB: data <= 32'hCFBEAE5D;	14'h10FC: data <= 32'hCFDC2C0F;	14'h10FD: data <= 32'hCFF9A9C2;	14'h10FE: data <= 32'hD0172774;	14'h10FF: data <= 32'hD034A527;	14'h1100: data <= 32'hD05222D9;	14'h1101: data <= 32'hD06FA08C;	14'h1102: data <= 32'hD08D1E3F;	14'h1103: data <= 32'hD0AA9BF1;	14'h1104: data <= 32'hD0C819A4;	14'h1105: data <= 32'hD0E59756;	14'h1106: data <= 32'hD1031509;	14'h1107: data <= 32'hD12092BB;	14'h1108: data <= 32'hD13E106E;	14'h1109: data <= 32'hD15B8E20;	14'h110A: data <= 32'hD1790BD3;	14'h110B: data <= 32'hD1968985;	14'h110C: data <= 32'hD1B39B66;	14'h110D: data <= 32'hD1CFF09A;	14'h110E: data <= 32'hD1EC45CD;	14'h110F: data <= 32'hD2089B00;	14'h1110: data <= 32'hD224F033;	14'h1111: data <= 32'hD2414567;	14'h1112: data <= 32'hD25D9A9A;	14'h1113: data <= 32'hD279EFCD;	14'h1114: data <= 32'hD2964500;	14'h1115: data <= 32'hD2B29A33;	14'h1116: data <= 32'hD2CEEF67;	14'h1117: data <= 32'hD2EB449A;	14'h1118: data <= 32'hD30799CD;	14'h1119: data <= 32'hD323EF00;	14'h111A: data <= 32'hD3404434;	14'h111B: data <= 32'hD35C9967;	14'h111C: data <= 32'hD378EE9A;	14'h111D: data <= 32'hD39543CD;	14'h111E: data <= 32'hD3B19900;	14'h111F: data <= 32'hD3CDEE34;	14'h1120: data <= 32'hD3EA4367;	14'h1121: data <= 32'hD406989A;	14'h1122: data <= 32'hD422EDCD;	14'h1123: data <= 32'hD43F4300;	14'h1124: data <= 32'hD45B9834;	14'h1125: data <= 32'hD477ED67;	14'h1126: data <= 32'hD494429A;	14'h1127: data <= 32'hD4B097CD;	14'h1128: data <= 32'hD4CCED01;	14'h1129: data <= 32'hD4E94234;	14'h112A: data <= 32'hD5058BC1;	14'h112B: data <= 32'hD52120C8;	14'h112C: data <= 32'hD53CB5CF;	14'h112D: data <= 32'hD5584AD5;	14'h112E: data <= 32'hD573DFDC;	14'h112F: data <= 32'hD58F74E2;	14'h1130: data <= 32'hD5AB09E9;	14'h1131: data <= 32'hD5C69EF0;	14'h1132: data <= 32'hD5E233F6;	14'h1133: data <= 32'hD5FDC8FD;	14'h1134: data <= 32'hD6195E04;	14'h1135: data <= 32'hD634F30A;	14'h1136: data <= 32'hD6508811;	14'h1137: data <= 32'hD66C1D17;	14'h1138: data <= 32'hD687B21E;	14'h1139: data <= 32'hD6A34725;	14'h113A: data <= 32'hD6BEDC2B;	14'h113B: data <= 32'hD6DA7132;	14'h113C: data <= 32'hD6F60639;	14'h113D: data <= 32'hD7119B3F;	14'h113E: data <= 32'hD72D3046;	14'h113F: data <= 32'hD748C54C;	14'h1140: data <= 32'hD7645A53;	14'h1141: data <= 32'hD77FEF5A;	14'h1142: data <= 32'hD79B8460;	14'h1143: data <= 32'hD7B71967;	14'h1144: data <= 32'hD7D2AE6D;	14'h1145: data <= 32'hD7EE4374;	14'h1146: data <= 32'hD809D87B;	14'h1147: data <= 32'hD8256D81;	14'h1148: data <= 32'hD8410288;	14'h1149: data <= 32'hD85D0C07;	14'h114A: data <= 32'hD8793ACB;	14'h114B: data <= 32'hD895698F;	14'h114C: data <= 32'hD8B19853;	14'h114D: data <= 32'hD8CDC716;	14'h114E: data <= 32'hD8E9F5DA;	14'h114F: data <= 32'hD906249E;	14'h1150: data <= 32'hD9225362;	14'h1151: data <= 32'hD93E8226;	14'h1152: data <= 32'hD95AB0EA;	14'h1153: data <= 32'hD976DFAE;	14'h1154: data <= 32'hD9930E72;	14'h1155: data <= 32'hD9AF3D36;	14'h1156: data <= 32'hD9CB6BFA;	14'h1157: data <= 32'hD9E79ABE;	14'h1158: data <= 32'hDA03C982;	14'h1159: data <= 32'hDA1FF846;	14'h115A: data <= 32'hDA3C270A;	14'h115B: data <= 32'hDA5855CE;	14'h115C: data <= 32'hDA748492;	14'h115D: data <= 32'hDA90B355;	14'h115E: data <= 32'hDAACE219;	14'h115F: data <= 32'hDAC910DD;	14'h1160: data <= 32'hDAE53FA1;	14'h1161: data <= 32'hDB016E65;	14'h1162: data <= 32'hDB1D9D29;	14'h1163: data <= 32'hDB39CBED;	14'h1164: data <= 32'hDB55FAB1;	14'h1165: data <= 32'hDB722975;	14'h1166: data <= 32'hDB8E5839;	14'h1167: data <= 32'hDBABD56C;	14'h1168: data <= 32'hDBCAE3F0;	14'h1169: data <= 32'hDBE9F275;	14'h116A: data <= 32'hDC0900F9;	14'h116B: data <= 32'hDC280F7E;	14'h116C: data <= 32'hDC471E02;	14'h116D: data <= 32'hDC662C87;	14'h116E: data <= 32'hDC853B0B;	14'h116F: data <= 32'hDCA44990;	14'h1170: data <= 32'hDCC35814;	14'h1171: data <= 32'hDCE26698;	14'h1172: data <= 32'hDD01751D;	14'h1173: data <= 32'hDD2083A1;	14'h1174: data <= 32'hDD3F9226;	14'h1175: data <= 32'hDD5EA0AA;	14'h1176: data <= 32'hDD7DAF2F;	14'h1177: data <= 32'hDD9CBDB3;	14'h1178: data <= 32'hDDBBCC38;	14'h1179: data <= 32'hDDDADABC;	14'h117A: data <= 32'hDDF9E941;	14'h117B: data <= 32'hDE18F7C5;	14'h117C: data <= 32'hDE38064A;	14'h117D: data <= 32'hDE5714CE;	14'h117E: data <= 32'hDE762353;	14'h117F: data <= 32'hDE9531D7;	14'h1180: data <= 32'hDEB4405C;	14'h1181: data <= 32'hDED34EE0;	14'h1182: data <= 32'hDEF25D65;	14'h1183: data <= 32'hDF116BE9;	14'h1184: data <= 32'hDF307A6E;	14'h1185: data <= 32'hDF505818;	14'h1186: data <= 32'hDF74BDCB;	14'h1187: data <= 32'hDF99237E;	14'h1188: data <= 32'hDFBD8931;	14'h1189: data <= 32'hDFE1EEE4;	14'h118A: data <= 32'hE0065497;	14'h118B: data <= 32'hE02ABA4A;	14'h118C: data <= 32'hE04F1FFD;	14'h118D: data <= 32'hE07385B0;	14'h118E: data <= 32'hE097EB63;	14'h118F: data <= 32'hE0BC5116;	14'h1190: data <= 32'hE0E0B6C9;	14'h1191: data <= 32'hE1051C7C;	14'h1192: data <= 32'hE129822F;	14'h1193: data <= 32'hE14DE7E2;	14'h1194: data <= 32'hE1724D95;	14'h1195: data <= 32'hE196B348;	14'h1196: data <= 32'hE1BB18FB;	14'h1197: data <= 32'hE1DF7EAE;	14'h1198: data <= 32'hE203E461;	14'h1199: data <= 32'hE2284A14;	14'h119A: data <= 32'hE24CAFC7;	14'h119B: data <= 32'hE271157A;	14'h119C: data <= 32'hE2957B2D;	14'h119D: data <= 32'hE2B9E0E0;	14'h119E: data <= 32'hE2DE4693;	14'h119F: data <= 32'hE302AC46;	14'h11A0: data <= 32'hE32711F9;	14'h11A1: data <= 32'hE34B77AC;	14'h11A2: data <= 32'hE36FDD5F;	14'h11A3: data <= 32'hE3944312;	14'h11A4: data <= 32'hE3BED417;	14'h11A5: data <= 32'hE3EA7F22;	14'h11A6: data <= 32'hE4162A2D;	14'h11A7: data <= 32'hE441D538;	14'h11A8: data <= 32'hE46D8043;	14'h11A9: data <= 32'hE4992B4E;	14'h11AA: data <= 32'hE4C4D659;	14'h11AB: data <= 32'hE4F08163;	14'h11AC: data <= 32'hE51C2C6E;	14'h11AD: data <= 32'hE547D779;	14'h11AE: data <= 32'hE5738284;	14'h11AF: data <= 32'hE59F2D8F;	14'h11B0: data <= 32'hE5CAD89A;	14'h11B1: data <= 32'hE5F683A5;	14'h11B2: data <= 32'hE6222EB0;	14'h11B3: data <= 32'hE64DD9BB;	14'h11B4: data <= 32'hE67984C6;	14'h11B5: data <= 32'hE6A52FD1;	14'h11B6: data <= 32'hE6D0DADB;	14'h11B7: data <= 32'hE6FC85E6;	14'h11B8: data <= 32'hE72830F1;	14'h11B9: data <= 32'hE753DBFC;	14'h11BA: data <= 32'hE77F8707;	14'h11BB: data <= 32'hE7AB3212;	14'h11BC: data <= 32'hE7D6DD1D;	14'h11BD: data <= 32'hE8028828;	14'h11BE: data <= 32'hE82E3333;	14'h11BF: data <= 32'hE859DE3E;	14'h11C0: data <= 32'hE8858949;	14'h11C1: data <= 32'hE8B13453;	14'h11C2: data <= 32'hE8E1BD42;	14'h11C3: data <= 32'hE916546D;	14'h11C4: data <= 32'hE94AEB98;	14'h11C5: data <= 32'hE97F82C4;	14'h11C6: data <= 32'hE9B419EF;	14'h11C7: data <= 32'hE9E8B11A;	14'h11C8: data <= 32'hEA1D4846;	14'h11C9: data <= 32'hEA51DF71;	14'h11CA: data <= 32'hEA86769C;	14'h11CB: data <= 32'hEABB0DC8;	14'h11CC: data <= 32'hEAEFA4F3;	14'h11CD: data <= 32'hEB243C1E;	14'h11CE: data <= 32'hEB58D34A;	14'h11CF: data <= 32'hEB8D6A75;	14'h11D0: data <= 32'hEBC201A0;	14'h11D1: data <= 32'hEBF698CC;	14'h11D2: data <= 32'hEC2B2FF7;	14'h11D3: data <= 32'hEC5FC722;	14'h11D4: data <= 32'hEC945E4E;	14'h11D5: data <= 32'hECC8F579;	14'h11D6: data <= 32'hECFD8CA4;	14'h11D7: data <= 32'hED3223D0;	14'h11D8: data <= 32'hED66BAFB;	14'h11D9: data <= 32'hED9B5227;	14'h11DA: data <= 32'hEDCFE952;	14'h11DB: data <= 32'hEE04807D;	14'h11DC: data <= 32'hEE3917A9;	14'h11DD: data <= 32'hEE6DAED4;	14'h11DE: data <= 32'hEEA245FF;	14'h11DF: data <= 32'hEED6DD2B;	14'h11E0: data <= 32'hEF0DE89B;	14'h11E1: data <= 32'hEF4C9F61;	14'h11E2: data <= 32'hEF8B5627;	14'h11E3: data <= 32'hEFCA0CED;	14'h11E4: data <= 32'hF008C3B3;	14'h11E5: data <= 32'hF0477A7A;	14'h11E6: data <= 32'hF0863140;	14'h11E7: data <= 32'hF0C4E806;	14'h11E8: data <= 32'hF1039ECC;	14'h11E9: data <= 32'hF1425593;	14'h11EA: data <= 32'hF1810C59;	14'h11EB: data <= 32'hF1BFC31F;	14'h11EC: data <= 32'hF1FE79E5;	14'h11ED: data <= 32'hF23D30AB;	14'h11EE: data <= 32'hF27BE772;	14'h11EF: data <= 32'hF2BA9E38;	14'h11F0: data <= 32'hF2F954FE;	14'h11F1: data <= 32'hF3380BC4;	14'h11F2: data <= 32'hF376C28B;	14'h11F3: data <= 32'hF3B57951;	14'h11F4: data <= 32'hF3F43017;	14'h11F5: data <= 32'hF432E6DD;	14'h11F6: data <= 32'hF4719DA3;	14'h11F7: data <= 32'hF4B0546A;	14'h11F8: data <= 32'hF4EF0B30;	14'h11F9: data <= 32'hF52DC1F6;	14'h11FA: data <= 32'hF56C78BC;	14'h11FB: data <= 32'hF5AB2F83;	14'h11FC: data <= 32'hF5E9E649;	14'h11FD: data <= 32'hF6289D0F;	14'h11FE: data <= 32'hF66753D5;	14'h11FF: data <= 32'hF6AFAC18;	14'h1200: data <= 32'hF6F8A36B;	14'h1201: data <= 32'hF7419ABE;	14'h1202: data <= 32'hF78A9211;	14'h1203: data <= 32'hF7D38964;	14'h1204: data <= 32'hF81C80B6;	14'h1205: data <= 32'hF8657809;	14'h1206: data <= 32'hF8AE6F5C;	14'h1207: data <= 32'hF8F766AF;	14'h1208: data <= 32'hF9405E02;	14'h1209: data <= 32'hF9895555;	14'h120A: data <= 32'hF9D24CA8;	14'h120B: data <= 32'hFA1B43FB;	14'h120C: data <= 32'hFA643B4E;	14'h120D: data <= 32'hFAAD32A1;	14'h120E: data <= 32'hFAF629F4;	14'h120F: data <= 32'hFB3F2146;	14'h1210: data <= 32'hFB881899;	14'h1211: data <= 32'hFBD10FEC;	14'h1212: data <= 32'hFC1A073F;	14'h1213: data <= 32'hFC62FE92;	14'h1214: data <= 32'hFCABF5E5;	14'h1215: data <= 32'hFCF4ED38;	14'h1216: data <= 32'hFD3DE48B;	14'h1217: data <= 32'hFD86DBDE;	14'h1218: data <= 32'hFDCFD331;	14'h1219: data <= 32'hFE18CA84;	14'h121A: data <= 32'hFE61C1D6;	14'h121B: data <= 32'hFEAAB929;	14'h121C: data <= 32'hFEF3B07C;	14'h121D: data <= 32'hFF426A4F;	14'h121E: data <= 32'hFF946EB4;	14'h121F: data <= 32'hFFE67319;	14'h1220: data <= 32'h0038777D;	14'h1221: data <= 32'h008A7BE2;	14'h1222: data <= 32'h00DC8047;	14'h1223: data <= 32'h012E84AC;	14'h1224: data <= 32'h01808910;	14'h1225: data <= 32'h01D28D75;	14'h1226: data <= 32'h022491DA;	14'h1227: data <= 32'h0276963F;	14'h1228: data <= 32'h02C89AA4;	14'h1229: data <= 32'h031A9F09;	14'h122A: data <= 32'h036CA36E;	14'h122B: data <= 32'h03BEA7D3;	14'h122C: data <= 32'h0410AC38;	14'h122D: data <= 32'h0462B09D;	14'h122E: data <= 32'h04B4B502;	14'h122F: data <= 32'h0506B967;	14'h1230: data <= 32'h0558BDCC;	14'h1231: data <= 32'h05AAC231;	14'h1232: data <= 32'h05FCC695;	14'h1233: data <= 32'h064ECAFA;	14'h1234: data <= 32'h06A0CF5F;	14'h1235: data <= 32'h06F2D3C4;	14'h1236: data <= 32'h0744D829;	14'h1237: data <= 32'h0796DC8E;	14'h1238: data <= 32'h07E8E0F3;	14'h1239: data <= 32'h083AE558;	14'h123A: data <= 32'h088CE9BD;	14'h123B: data <= 32'h08E16B0D;	14'h123C: data <= 32'h093AE635;	14'h123D: data <= 32'h0994615C;	14'h123E: data <= 32'h09EDDC84;	14'h123F: data <= 32'h0A4757AB;	14'h1240: data <= 32'h0AA0D2D3;	14'h1241: data <= 32'h0AFA4DFA;	14'h1242: data <= 32'h0B53C922;	14'h1243: data <= 32'h0BAD4449;	14'h1244: data <= 32'h0C06BF71;	14'h1245: data <= 32'h0C603A98;	14'h1246: data <= 32'h0CB9B5C0;	14'h1247: data <= 32'h0D1330E7;	14'h1248: data <= 32'h0D6CAC0F;	14'h1249: data <= 32'h0DC62736;	14'h124A: data <= 32'h0E1FA25E;	14'h124B: data <= 32'h0E791D85;	14'h124C: data <= 32'h0ED298AD;	14'h124D: data <= 32'h0F2C13D4;	14'h124E: data <= 32'h0F858EFC;	14'h124F: data <= 32'h0FDF0A23;	14'h1250: data <= 32'h1038854B;	14'h1251: data <= 32'h10920072;	14'h1252: data <= 32'h10EB7B9A;	14'h1253: data <= 32'h1144F6C1;	14'h1254: data <= 32'h119E71E9;	14'h1255: data <= 32'h11F7ED10;	14'h1256: data <= 32'h12516838;	14'h1257: data <= 32'h12AAE35F;	14'h1258: data <= 32'h13045E87;	14'h1259: data <= 32'h135E0148;	14'h125A: data <= 32'h13BC9738;	14'h125B: data <= 32'h141B2D28;	14'h125C: data <= 32'h1479C318;	14'h125D: data <= 32'h14D85909;	14'h125E: data <= 32'h1536EEF9;	14'h125F: data <= 32'h159584E9;	14'h1260: data <= 32'h15F41AD9;	14'h1261: data <= 32'h1652B0C9;	14'h1262: data <= 32'h16B146B9;	14'h1263: data <= 32'h170FDCA9;	14'h1264: data <= 32'h176E729A;	14'h1265: data <= 32'h17CD088A;	14'h1266: data <= 32'h182B9E7A;	14'h1267: data <= 32'h188A346A;	14'h1268: data <= 32'h18E8CA5A;	14'h1269: data <= 32'h1947604A;	14'h126A: data <= 32'h19A5F63A;	14'h126B: data <= 32'h1A048C2B;	14'h126C: data <= 32'h1A63221B;	14'h126D: data <= 32'h1AC1B80B;	14'h126E: data <= 32'h1B204DFB;	14'h126F: data <= 32'h1B7EE3EB;	14'h1270: data <= 32'h1BDD79DB;	14'h1271: data <= 32'h1C3C0FCB;	14'h1272: data <= 32'h1C9AA5BC;	14'h1273: data <= 32'h1CF93BAC;	14'h1274: data <= 32'h1D57D19C;	14'h1275: data <= 32'h1DB6678C;	14'h1276: data <= 32'h1E14FD7C;	14'h1277: data <= 32'h1E73936C;	14'h1278: data <= 32'h1ED398BD;	14'h1279: data <= 32'h1F3427D2;	14'h127A: data <= 32'h1F94B6E7;	14'h127B: data <= 32'h1FF545FC;	14'h127C: data <= 32'h2055D511;	14'h127D: data <= 32'h20B66425;	14'h127E: data <= 32'h2116F33A;	14'h127F: data <= 32'h2177824F;	14'h1280: data <= 32'h21D81164;	14'h1281: data <= 32'h2238A079;	14'h1282: data <= 32'h22992F8E;	14'h1283: data <= 32'h22F9BEA3;	14'h1284: data <= 32'h235A4DB8;	14'h1285: data <= 32'h23BADCCD;	14'h1286: data <= 32'h241B6BE1;	14'h1287: data <= 32'h247BFAF6;	14'h1288: data <= 32'h24DC8A0B;	14'h1289: data <= 32'h253D1920;	14'h128A: data <= 32'h259DA835;	14'h128B: data <= 32'h25FE374A;	14'h128C: data <= 32'h265EC65F;	14'h128D: data <= 32'h26BF5574;	14'h128E: data <= 32'h271FE489;	14'h128F: data <= 32'h2780739D;	14'h1290: data <= 32'h27E102B2;	14'h1291: data <= 32'h284191C7;	14'h1292: data <= 32'h28A220DC;	14'h1293: data <= 32'h2902AFF1;	14'h1294: data <= 32'h29633F06;	14'h1295: data <= 32'h29C3CE1B;	14'h1296: data <= 32'h2A23C5C7;	14'h1297: data <= 32'h2A82EFF6;	14'h1298: data <= 32'h2AE21A26;	14'h1299: data <= 32'h2B414456;	14'h129A: data <= 32'h2BA06E86;	14'h129B: data <= 32'h2BFF98B6;	14'h129C: data <= 32'h2C5EC2E6;	14'h129D: data <= 32'h2CBDED15;	14'h129E: data <= 32'h2D1D1745;	14'h129F: data <= 32'h2D7C4175;	14'h12A0: data <= 32'h2DDB6BA5;	14'h12A1: data <= 32'h2E3A95D5;	14'h12A2: data <= 32'h2E99C005;	14'h12A3: data <= 32'h2EF8EA34;	14'h12A4: data <= 32'h2F581464;	14'h12A5: data <= 32'h2FB73E94;	14'h12A6: data <= 32'h301668C4;	14'h12A7: data <= 32'h307592F4;	14'h12A8: data <= 32'h30D4BD24;	14'h12A9: data <= 32'h3133E753;	14'h12AA: data <= 32'h31931183;	14'h12AB: data <= 32'h31F23BB3;	14'h12AC: data <= 32'h325165E3;	14'h12AD: data <= 32'h32B09013;	14'h12AE: data <= 32'h330FBA43;	14'h12AF: data <= 32'h336EE472;	14'h12B0: data <= 32'h33CE0EA2;	14'h12B1: data <= 32'h342D38D2;	14'h12B2: data <= 32'h348C6302;	14'h12B3: data <= 32'h34EB8D32;	14'h12B4: data <= 32'h354A4792;	14'h12B5: data <= 32'h35A5D752;	14'h12B6: data <= 32'h36016713;	14'h12B7: data <= 32'h365CF6D3;	14'h12B8: data <= 32'h36B88693;	14'h12B9: data <= 32'h37141654;	14'h12BA: data <= 32'h376FA614;	14'h12BB: data <= 32'h37CB35D4;	14'h12BC: data <= 32'h3826C594;	14'h12BD: data <= 32'h38825555;	14'h12BE: data <= 32'h38DDE515;	14'h12BF: data <= 32'h393974D5;	14'h12C0: data <= 32'h39950495;	14'h12C1: data <= 32'h39F09456;	14'h12C2: data <= 32'h3A4C2416;	14'h12C3: data <= 32'h3AA7B3D6;	14'h12C4: data <= 32'h3B034397;	14'h12C5: data <= 32'h3B5ED357;	14'h12C6: data <= 32'h3BBA6317;	14'h12C7: data <= 32'h3C15F2D7;	14'h12C8: data <= 32'h3C718298;	14'h12C9: data <= 32'h3CCD1258;	14'h12CA: data <= 32'h3D28A218;	14'h12CB: data <= 32'h3D8431D9;	14'h12CC: data <= 32'h3DDFC199;	14'h12CD: data <= 32'h3E3B5159;	14'h12CE: data <= 32'h3E96E119;	14'h12CF: data <= 32'h3EF270DA;	14'h12D0: data <= 32'h3F4E009A;	14'h12D1: data <= 32'h3FA9905A;	14'h12D2: data <= 32'h4005201B;	14'h12D3: data <= 32'h405C2454;	14'h12D4: data <= 32'h40B225FE;	14'h12D5: data <= 32'h410827A7;	14'h12D6: data <= 32'h415E2951;	14'h12D7: data <= 32'h41B42AFA;	14'h12D8: data <= 32'h420A2CA4;	14'h12D9: data <= 32'h42602E4E;	14'h12DA: data <= 32'h42B62FF7;	14'h12DB: data <= 32'h430C31A1;	14'h12DC: data <= 32'h4362334A;	14'h12DD: data <= 32'h43B834F4;	14'h12DE: data <= 32'h440E369E;	14'h12DF: data <= 32'h44643847;	14'h12E0: data <= 32'h44BA39F1;	14'h12E1: data <= 32'h45103B9A;	14'h12E2: data <= 32'h45663D44;	14'h12E3: data <= 32'h45BC3EEE;	14'h12E4: data <= 32'h46124097;	14'h12E5: data <= 32'h46684241;	14'h12E6: data <= 32'h46BE43EA;	14'h12E7: data <= 32'h47144594;	14'h12E8: data <= 32'h476A473E;	14'h12E9: data <= 32'h47C048E7;	14'h12EA: data <= 32'h48164A91;	14'h12EB: data <= 32'h486C4C3B;	14'h12EC: data <= 32'h48C24DE4;	14'h12ED: data <= 32'h49184F8E;	14'h12EE: data <= 32'h496E5137;	14'h12EF: data <= 32'h49C452E1;	14'h12F0: data <= 32'h4A1A548B;	14'h12F1: data <= 32'h4A6C509E;	14'h12F2: data <= 32'h4ABA83AB;	14'h12F3: data <= 32'h4B08B6B8;	14'h12F4: data <= 32'h4B56E9C6;	14'h12F5: data <= 32'h4BA51CD3;	14'h12F6: data <= 32'h4BF34FE0;	14'h12F7: data <= 32'h4C4182EE;	14'h12F8: data <= 32'h4C8FB5FB;	14'h12F9: data <= 32'h4CDDE908;	14'h12FA: data <= 32'h4D2C1C15;	14'h12FB: data <= 32'h4D7A4F23;	14'h12FC: data <= 32'h4DC88230;	14'h12FD: data <= 32'h4E16B53D;	14'h12FE: data <= 32'h4E64E84B;	14'h12FF: data <= 32'h4EB31B58;	14'h1300: data <= 32'h4F014E65;	14'h1301: data <= 32'h4F4F8173;	14'h1302: data <= 32'h4F9DB480;	14'h1303: data <= 32'h4FEBE78D;	14'h1304: data <= 32'h503A1A9A;	14'h1305: data <= 32'h50884DA8;	14'h1306: data <= 32'h50D680B5;	14'h1307: data <= 32'h5124B3C2;	14'h1308: data <= 32'h5172E6D0;	14'h1309: data <= 32'h51C119DD;	14'h130A: data <= 32'h520F4CEA;	14'h130B: data <= 32'h525D7FF8;	14'h130C: data <= 32'h52ABB305;	14'h130D: data <= 32'h52F9E612;	14'h130E: data <= 32'h5348191F;	14'h130F: data <= 32'h5394642B;	14'h1310: data <= 32'h53D99A9F;	14'h1311: data <= 32'h541ED113;	14'h1312: data <= 32'h54640787;	14'h1313: data <= 32'h54A93DFB;	14'h1314: data <= 32'h54EE746F;	14'h1315: data <= 32'h5533AAE3;	14'h1316: data <= 32'h5578E157;	14'h1317: data <= 32'h55BE17CB;	14'h1318: data <= 32'h56034E3F;	14'h1319: data <= 32'h564884B3;	14'h131A: data <= 32'h568DBB27;	14'h131B: data <= 32'h56D2F19B;	14'h131C: data <= 32'h5718280F;	14'h131D: data <= 32'h575D5E83;	14'h131E: data <= 32'h57A294F7;	14'h131F: data <= 32'h57E7CB6B;	14'h1320: data <= 32'h582D01DF;	14'h1321: data <= 32'h58723853;	14'h1322: data <= 32'h58B76EC7;	14'h1323: data <= 32'h58FCA53B;	14'h1324: data <= 32'h5941DBAF;	14'h1325: data <= 32'h59871223;	14'h1326: data <= 32'h59CC4897;	14'h1327: data <= 32'h5A117F0B;	14'h1328: data <= 32'h5A56B57F;	14'h1329: data <= 32'h5A9BEBF3;	14'h132A: data <= 32'h5AE12267;	14'h132B: data <= 32'h5B2658DB;	14'h132C: data <= 32'h5B6B8F4F;	14'h132D: data <= 32'h5BB0C5C3;	14'h132E: data <= 32'h5BEDF8B1;	14'h132F: data <= 32'h5C2A5E79;	14'h1330: data <= 32'h5C66C441;	14'h1331: data <= 32'h5CA32A08;	14'h1332: data <= 32'h5CDF8FD0;	14'h1333: data <= 32'h5D1BF598;	14'h1334: data <= 32'h5D585B60;	14'h1335: data <= 32'h5D94C127;	14'h1336: data <= 32'h5DD126EF;	14'h1337: data <= 32'h5E0D8CB7;	14'h1338: data <= 32'h5E49F27E;	14'h1339: data <= 32'h5E865846;	14'h133A: data <= 32'h5EC2BE0E;	14'h133B: data <= 32'h5EFF23D5;	14'h133C: data <= 32'h5F3B899D;	14'h133D: data <= 32'h5F77EF65;	14'h133E: data <= 32'h5FB4552C;	14'h133F: data <= 32'h5FF0BAF4;	14'h1340: data <= 32'h602D20BC;	14'h1341: data <= 32'h60698684;	14'h1342: data <= 32'h60A5EC4B;	14'h1343: data <= 32'h60E25213;	14'h1344: data <= 32'h611EB7DB;	14'h1345: data <= 32'h615B1DA2;	14'h1346: data <= 32'h6197836A;	14'h1347: data <= 32'h61D3E932;	14'h1348: data <= 32'h62104EF9;	14'h1349: data <= 32'h624CB4C1;	14'h134A: data <= 32'h62891A89;	14'h134B: data <= 32'h62C58050;	14'h134C: data <= 32'h62FD02E2;	14'h134D: data <= 32'h6331582A;	14'h134E: data <= 32'h6365AD72;	14'h134F: data <= 32'h639A02BA;	14'h1350: data <= 32'h63CE5802;	14'h1351: data <= 32'h6402AD4A;	14'h1352: data <= 32'h64370292;	14'h1353: data <= 32'h646B57DA;	14'h1354: data <= 32'h649FAD22;	14'h1355: data <= 32'h64D4026A;	14'h1356: data <= 32'h650857B2;	14'h1357: data <= 32'h653CACFA;	14'h1358: data <= 32'h65710241;	14'h1359: data <= 32'h65A55789;	14'h135A: data <= 32'h65D9ACD1;	14'h135B: data <= 32'h660E0219;	14'h135C: data <= 32'h66425761;	14'h135D: data <= 32'h6676ACA9;	14'h135E: data <= 32'h66AB01F1;	14'h135F: data <= 32'h66DF5739;	14'h1360: data <= 32'h6713AC81;	14'h1361: data <= 32'h674801C9;	14'h1362: data <= 32'h677C5711;	14'h1363: data <= 32'h67B0AC59;	14'h1364: data <= 32'h67E501A1;	14'h1365: data <= 32'h681956E9;	14'h1366: data <= 32'h684DAC31;	14'h1367: data <= 32'h68820179;	14'h1368: data <= 32'h68B656C1;	14'h1369: data <= 32'h68EAAC09;	14'h136A: data <= 32'h691CD741;	14'h136B: data <= 32'h694A0823;	14'h136C: data <= 32'h69773905;	14'h136D: data <= 32'h69A469E6;	14'h136E: data <= 32'h69D19AC8;	14'h136F: data <= 32'h69FECBAA;	14'h1370: data <= 32'h6A2BFC8B;	14'h1371: data <= 32'h6A592D6D;	14'h1372: data <= 32'h6A865E4F;	14'h1373: data <= 32'h6AB38F30;	14'h1374: data <= 32'h6AE0C012;	14'h1375: data <= 32'h6B0DF0F4;	14'h1376: data <= 32'h6B3B21D5;	14'h1377: data <= 32'h6B6852B7;	14'h1378: data <= 32'h6B958399;	14'h1379: data <= 32'h6BC2B47A;	14'h137A: data <= 32'h6BEFE55C;	14'h137B: data <= 32'h6C1D163E;	14'h137C: data <= 32'h6C4A471F;	14'h137D: data <= 32'h6C777801;	14'h137E: data <= 32'h6CA4A8E3;	14'h137F: data <= 32'h6CD1D9C4;	14'h1380: data <= 32'h6CFF0AA6;	14'h1381: data <= 32'h6D2C3B88;	14'h1382: data <= 32'h6D596C69;	14'h1383: data <= 32'h6D869D4B;	14'h1384: data <= 32'h6DB3CE2D;	14'h1385: data <= 32'h6DE0FF0E;	14'h1386: data <= 32'h6E0E2FF0;	14'h1387: data <= 32'h6E3B60D2;	14'h1388: data <= 32'h6E6891B4;	14'h1389: data <= 32'h6E8FBBB3;	14'h138A: data <= 32'h6EB6E5B2;	14'h138B: data <= 32'h6EDE0FB2;	14'h138C: data <= 32'h6F0539B1;	14'h138D: data <= 32'h6F2C63B1;	14'h138E: data <= 32'h6F538DB0;	14'h138F: data <= 32'h6F7AB7B0;	14'h1390: data <= 32'h6FA1E1AF;	14'h1391: data <= 32'h6FC90BAF;	14'h1392: data <= 32'h6FF035AE;	14'h1393: data <= 32'h70175FAE;	14'h1394: data <= 32'h703E89AD;	14'h1395: data <= 32'h7065B3AD;	14'h1396: data <= 32'h708CDDAC;	14'h1397: data <= 32'h70B407AC;	14'h1398: data <= 32'h70DB31AB;	14'h1399: data <= 32'h71025BAB;	14'h139A: data <= 32'h712985AA;	14'h139B: data <= 32'h7150AFAA;	14'h139C: data <= 32'h7177D9A9;	14'h139D: data <= 32'h719F03A9;	14'h139E: data <= 32'h71C62DA8;	14'h139F: data <= 32'h71ED57A8;	14'h13A0: data <= 32'h721481A7;	14'h13A1: data <= 32'h723BABA7;	14'h13A2: data <= 32'h7262D5A6;	14'h13A3: data <= 32'h7289FFA6;	14'h13A4: data <= 32'h72B129A5;	14'h13A5: data <= 32'h72D853A5;	14'h13A6: data <= 32'h72FF7DA4;	14'h13A7: data <= 32'h7322CC50;	14'h13A8: data <= 32'h73446DB7;	14'h13A9: data <= 32'h73660F1D;	14'h13AA: data <= 32'h7387B084;	14'h13AB: data <= 32'h73A951EA;	14'h13AC: data <= 32'h73CAF351;	14'h13AD: data <= 32'h73EC94B7;	14'h13AE: data <= 32'h740E361E;	14'h13AF: data <= 32'h742FD784;	14'h13B0: data <= 32'h745178EA;	14'h13B1: data <= 32'h74731A51;	14'h13B2: data <= 32'h7494BBB7;	14'h13B3: data <= 32'h74B65D1E;	14'h13B4: data <= 32'h74D7FE84;	14'h13B5: data <= 32'h74F99FEB;	14'h13B6: data <= 32'h751B4151;	14'h13B7: data <= 32'h753CE2B8;	14'h13B8: data <= 32'h755E841E;	14'h13B9: data <= 32'h75802585;	14'h13BA: data <= 32'h75A1C6EB;	14'h13BB: data <= 32'h75C36852;	14'h13BC: data <= 32'h75E509B8;	14'h13BD: data <= 32'h7606AB1F;	14'h13BE: data <= 32'h76284C85;	14'h13BF: data <= 32'h7649EDEC;	14'h13C0: data <= 32'h766B8F52;	14'h13C1: data <= 32'h768D30B9;	14'h13C2: data <= 32'h76AED21F;	14'h13C3: data <= 32'h76D07386;	14'h13C4: data <= 32'h76F214EC;	14'h13C5: data <= 32'h771176F7;	14'h13C6: data <= 32'h772D63D7;	14'h13C7: data <= 32'h774950B8;	14'h13C8: data <= 32'h77653D98;	14'h13C9: data <= 32'h77812A79;	14'h13CA: data <= 32'h779D1759;	14'h13CB: data <= 32'h77B9043A;	14'h13CC: data <= 32'h77D4F11A;	14'h13CD: data <= 32'h77F0DDFB;	14'h13CE: data <= 32'h780CCADB;	14'h13CF: data <= 32'h7828B7BC;	14'h13D0: data <= 32'h7844A49C;	14'h13D1: data <= 32'h7860917D;	14'h13D2: data <= 32'h787C7E5D;	14'h13D3: data <= 32'h78986B3E;	14'h13D4: data <= 32'h78B4581E;	14'h13D5: data <= 32'h78D044FF;	14'h13D6: data <= 32'h78EC31DF;	14'h13D7: data <= 32'h79081EC0;	14'h13D8: data <= 32'h79240BA0;	14'h13D9: data <= 32'h793FF881;	14'h13DA: data <= 32'h795BE561;	14'h13DB: data <= 32'h7977D242;	14'h13DC: data <= 32'h7993BF22;	14'h13DD: data <= 32'h79AFAC02;	14'h13DE: data <= 32'h79CB98E3;	14'h13DF: data <= 32'h79E785C3;	14'h13E0: data <= 32'h7A0372A4;	14'h13E1: data <= 32'h7A1F5F84;	14'h13E2: data <= 32'h7A3B4C65;	14'h13E3: data <= 32'h7A56B280;	14'h13E4: data <= 32'h7A6CD4E4;	14'h13E5: data <= 32'h7A82F748;	14'h13E6: data <= 32'h7A9919AC;	14'h13E7: data <= 32'h7AAF3C10;	14'h13E8: data <= 32'h7AC55E74;	14'h13E9: data <= 32'h7ADB80D9;	14'h13EA: data <= 32'h7AF1A33D;	14'h13EB: data <= 32'h7B07C5A1;	14'h13EC: data <= 32'h7B1DE805;	14'h13ED: data <= 32'h7B340A69;	14'h13EE: data <= 32'h7B4A2CCD;	14'h13EF: data <= 32'h7B604F31;	14'h13F0: data <= 32'h7B767195;	14'h13F1: data <= 32'h7B8C93F9;	14'h13F2: data <= 32'h7BA2B65E;	14'h13F3: data <= 32'h7BB8D8C2;	14'h13F4: data <= 32'h7BCEFB26;	14'h13F5: data <= 32'h7BE51D8A;	14'h13F6: data <= 32'h7BFB3FEE;	14'h13F7: data <= 32'h7C116252;	14'h13F8: data <= 32'h7C2784B6;	14'h13F9: data <= 32'h7C3DA71A;	14'h13FA: data <= 32'h7C53C97E;	14'h13FB: data <= 32'h7C69EBE3;	14'h13FC: data <= 32'h7C800E47;	14'h13FD: data <= 32'h7C9630AB;	14'h13FE: data <= 32'h7CAC530F;	14'h13FF: data <= 32'h7CC27573;	14'h1400: data <= 32'h7CD897D7;	14'h1401: data <= 32'h7CEEBA3B;	14'h1402: data <= 32'h7D002158;	14'h1403: data <= 32'h7D104257;	14'h1404: data <= 32'h7D206357;	14'h1405: data <= 32'h7D308456;	14'h1406: data <= 32'h7D40A556;	14'h1407: data <= 32'h7D50C655;	14'h1408: data <= 32'h7D60E755;	14'h1409: data <= 32'h7D710854;	14'h140A: data <= 32'h7D812954;	14'h140B: data <= 32'h7D914A53;	14'h140C: data <= 32'h7DA16B53;	14'h140D: data <= 32'h7DB18C52;	14'h140E: data <= 32'h7DC1AD52;	14'h140F: data <= 32'h7DD1CE51;	14'h1410: data <= 32'h7DE1EF51;	14'h1411: data <= 32'h7DF21050;	14'h1412: data <= 32'h7E023150;	14'h1413: data <= 32'h7E12524F;	14'h1414: data <= 32'h7E22734F;	14'h1415: data <= 32'h7E32944E;	14'h1416: data <= 32'h7E42B54E;	14'h1417: data <= 32'h7E52D64D;	14'h1418: data <= 32'h7E62F74D;	14'h1419: data <= 32'h7E73184C;	14'h141A: data <= 32'h7E83394C;	14'h141B: data <= 32'h7E935A4B;	14'h141C: data <= 32'h7EA37B4B;	14'h141D: data <= 32'h7EB39C4A;	14'h141E: data <= 32'h7EC3BD4A;	14'h141F: data <= 32'h7ED3DE49;	14'h1420: data <= 32'h7EE09E16;	14'h1421: data <= 32'h7EE9C69C;	14'h1422: data <= 32'h7EF2EF22;	14'h1423: data <= 32'h7EFC17A8;	14'h1424: data <= 32'h7F05402E;	14'h1425: data <= 32'h7F0E68B5;	14'h1426: data <= 32'h7F17913B;	14'h1427: data <= 32'h7F20B9C1;	14'h1428: data <= 32'h7F29E247;	14'h1429: data <= 32'h7F330ACD;	14'h142A: data <= 32'h7F3C3354;	14'h142B: data <= 32'h7F455BDA;	14'h142C: data <= 32'h7F4E8460;	14'h142D: data <= 32'h7F57ACE6;	14'h142E: data <= 32'h7F60D56C;	14'h142F: data <= 32'h7F69FDF3;	14'h1430: data <= 32'h7F732679;	14'h1431: data <= 32'h7F7C4EFF;	14'h1432: data <= 32'h7F857785;	14'h1433: data <= 32'h7F8EA00B;	14'h1434: data <= 32'h7F97C892;	14'h1435: data <= 32'h7FA0F118;	14'h1436: data <= 32'h7FAA199E;	14'h1437: data <= 32'h7FB34224;	14'h1438: data <= 32'h7FBC6AAA;	14'h1439: data <= 32'h7FC59330;	14'h143A: data <= 32'h7FCEBBB7;	14'h143B: data <= 32'h7FD7E43D;	14'h143C: data <= 32'h7FE10CC3;	14'h143D: data <= 32'h7FEA3549;	14'h143E: data <= 32'h7FF1C97F;	14'h143F: data <= 32'h7FF2424B;	14'h1440: data <= 32'h7FF2BB16;	14'h1441: data <= 32'h7FF333E2;	14'h1442: data <= 32'h7FF3ACAD;	14'h1443: data <= 32'h7FF42579;	14'h1444: data <= 32'h7FF49E44;	14'h1445: data <= 32'h7FF51710;	14'h1446: data <= 32'h7FF58FDC;	14'h1447: data <= 32'h7FF608A7;	14'h1448: data <= 32'h7FF68173;	14'h1449: data <= 32'h7FF6FA3E;	14'h144A: data <= 32'h7FF7730A;	14'h144B: data <= 32'h7FF7EBD5;	14'h144C: data <= 32'h7FF864A1;	14'h144D: data <= 32'h7FF8DD6D;	14'h144E: data <= 32'h7FF95638;	14'h144F: data <= 32'h7FF9CF04;	14'h1450: data <= 32'h7FFA47CF;	14'h1451: data <= 32'h7FFAC09B;	14'h1452: data <= 32'h7FFB3966;	14'h1453: data <= 32'h7FFBB232;	14'h1454: data <= 32'h7FFC2AFE;	14'h1455: data <= 32'h7FFCA3C9;	14'h1456: data <= 32'h7FFD1C95;	14'h1457: data <= 32'h7FFD9560;	14'h1458: data <= 32'h7FFE0E2C;	14'h1459: data <= 32'h7FFE86F7;	14'h145A: data <= 32'h7FFEFFC3;	14'h145B: data <= 32'h7FFF788F;	14'h145C: data <= 32'h7FFFF15A;	14'h145D: data <= 32'h7FF72900;	14'h145E: data <= 32'h7FED19DD;	14'h145F: data <= 32'h7FE30ABB;	14'h1460: data <= 32'h7FD8FB99;	14'h1461: data <= 32'h7FCEEC77;	14'h1462: data <= 32'h7FC4DD55;	14'h1463: data <= 32'h7FBACE33;	14'h1464: data <= 32'h7FB0BF11;	14'h1465: data <= 32'h7FA6AFEF;	14'h1466: data <= 32'h7F9CA0CD;	14'h1467: data <= 32'h7F9291AB;	14'h1468: data <= 32'h7F888288;	14'h1469: data <= 32'h7F7E7366;	14'h146A: data <= 32'h7F746444;	14'h146B: data <= 32'h7F6A5522;	14'h146C: data <= 32'h7F604600;	14'h146D: data <= 32'h7F5636DE;	14'h146E: data <= 32'h7F4C27BC;	14'h146F: data <= 32'h7F42189A;	14'h1470: data <= 32'h7F380978;	14'h1471: data <= 32'h7F2DFA56;	14'h1472: data <= 32'h7F23EB33;	14'h1473: data <= 32'h7F19DC11;	14'h1474: data <= 32'h7F0FCCEF;	14'h1475: data <= 32'h7F05BDCD;	14'h1476: data <= 32'h7EFBAEAB;	14'h1477: data <= 32'h7EF19F89;	14'h1478: data <= 32'h7EE79067;	14'h1479: data <= 32'h7EDD8145;	14'h147A: data <= 32'h7ED37223;	14'h147B: data <= 32'h7EC25C38;	14'h147C: data <= 32'h7EAC18E2;	14'h147D: data <= 32'h7E95D58C;	14'h147E: data <= 32'h7E7F9237;	14'h147F: data <= 32'h7E694EE1;	14'h1480: data <= 32'h7E530B8B;	14'h1481: data <= 32'h7E3CC835;	14'h1482: data <= 32'h7E2684E0;	14'h1483: data <= 32'h7E10418A;	14'h1484: data <= 32'h7DF9FE34;	14'h1485: data <= 32'h7DE3BADE;	14'h1486: data <= 32'h7DCD7788;	14'h1487: data <= 32'h7DB73433;	14'h1488: data <= 32'h7DA0F0DD;	14'h1489: data <= 32'h7D8AAD87;	14'h148A: data <= 32'h7D746A31;	14'h148B: data <= 32'h7D5E26DB;	14'h148C: data <= 32'h7D47E386;	14'h148D: data <= 32'h7D31A030;	14'h148E: data <= 32'h7D1B5CDA;	14'h148F: data <= 32'h7D051984;	14'h1490: data <= 32'h7CEED62E;	14'h1491: data <= 32'h7CD892D9;	14'h1492: data <= 32'h7CC24F83;	14'h1493: data <= 32'h7CAC0C2D;	14'h1494: data <= 32'h7C95C8D7;	14'h1495: data <= 32'h7C7F8581;	14'h1496: data <= 32'h7C69422C;	14'h1497: data <= 32'h7C52FED6;	14'h1498: data <= 32'h7C3CBB80;	14'h1499: data <= 32'h7C22C2C6;	14'h149A: data <= 32'h7BFEE658;	14'h149B: data <= 32'h7BDB09E9;	14'h149C: data <= 32'h7BB72D7B;	14'h149D: data <= 32'h7B93510C;	14'h149E: data <= 32'h7B6F749E;	14'h149F: data <= 32'h7B4B982F;	14'h14A0: data <= 32'h7B27BBC1;	14'h14A1: data <= 32'h7B03DF52;	14'h14A2: data <= 32'h7AE002E4;	14'h14A3: data <= 32'h7ABC2675;	14'h14A4: data <= 32'h7A984A07;	14'h14A5: data <= 32'h7A746D98;	14'h14A6: data <= 32'h7A509129;	14'h14A7: data <= 32'h7A2CB4BB;	14'h14A8: data <= 32'h7A08D84C;	14'h14A9: data <= 32'h79E4FBDE;	14'h14AA: data <= 32'h79C11F6F;	14'h14AB: data <= 32'h799D4301;	14'h14AC: data <= 32'h79796692;	14'h14AD: data <= 32'h79558A24;	14'h14AE: data <= 32'h7931ADB5;	14'h14AF: data <= 32'h790DD147;	14'h14B0: data <= 32'h78E9F4D8;	14'h14B1: data <= 32'h78C6186A;	14'h14B2: data <= 32'h78A23BFB;	14'h14B3: data <= 32'h787E5F8D;	14'h14B4: data <= 32'h785A831E;	14'h14B5: data <= 32'h7836A6AF;	14'h14B6: data <= 32'h7812CA41;	14'h14B7: data <= 32'h77EEEDD2;	14'h14B8: data <= 32'h77BDAC8A;	14'h14B9: data <= 32'h778C001A;	14'h14BA: data <= 32'h775A53AB;	14'h14BB: data <= 32'h7728A73B;	14'h14BC: data <= 32'h76F6FACC;	14'h14BD: data <= 32'h76C54E5C;	14'h14BE: data <= 32'h7693A1ED;	14'h14BF: data <= 32'h7661F57D;	14'h14C0: data <= 32'h7630490D;	14'h14C1: data <= 32'h75FE9C9E;	14'h14C2: data <= 32'h75CCF02E;	14'h14C3: data <= 32'h759B43BF;	14'h14C4: data <= 32'h7569974F;	14'h14C5: data <= 32'h7537EAE0;	14'h14C6: data <= 32'h75063E70;	14'h14C7: data <= 32'h74D49201;	14'h14C8: data <= 32'h74A2E591;	14'h14C9: data <= 32'h74713922;	14'h14CA: data <= 32'h743F8CB2;	14'h14CB: data <= 32'h740DE043;	14'h14CC: data <= 32'h73DC33D3;	14'h14CD: data <= 32'h73AA8764;	14'h14CE: data <= 32'h7378DAF4;	14'h14CF: data <= 32'h73472E85;	14'h14D0: data <= 32'h73158215;	14'h14D1: data <= 32'h72E3D5A5;	14'h14D2: data <= 32'h72B22936;	14'h14D3: data <= 32'h72807CC6;	14'h14D4: data <= 32'h724ED057;	14'h14D5: data <= 32'h721D23E7;	14'h14D6: data <= 32'h71E2C992;	14'h14D7: data <= 32'h71A41849;	14'h14D8: data <= 32'h71656701;	14'h14D9: data <= 32'h7126B5B8;	14'h14DA: data <= 32'h70E8046F;	14'h14DB: data <= 32'h70A95327;	14'h14DC: data <= 32'h706AA1DE;	14'h14DD: data <= 32'h702BF095;	14'h14DE: data <= 32'h6FED3F4D;	14'h14DF: data <= 32'h6FAE8E04;	14'h14E0: data <= 32'h6F6FDCBC;	14'h14E1: data <= 32'h6F312B73;	14'h14E2: data <= 32'h6EF27A2A;	14'h14E3: data <= 32'h6EB3C8E2;	14'h14E4: data <= 32'h6E751799;	14'h14E5: data <= 32'h6E366650;	14'h14E6: data <= 32'h6DF7B508;	14'h14E7: data <= 32'h6DB903BF;	14'h14E8: data <= 32'h6D7A5277;	14'h14E9: data <= 32'h6D3BA12E;	14'h14EA: data <= 32'h6CFCEFE5;	14'h14EB: data <= 32'h6CBE3E9D;	14'h14EC: data <= 32'h6C7F8D54;	14'h14ED: data <= 32'h6C40DC0B;	14'h14EE: data <= 32'h6C022AC3;	14'h14EF: data <= 32'h6BC3797A;	14'h14F0: data <= 32'h6B84C832;	14'h14F1: data <= 32'h6B4616E9;	14'h14F2: data <= 32'h6B0765A0;	14'h14F3: data <= 32'h6AC8B458;	14'h14F4: data <= 32'h6A85DEDB;	14'h14F5: data <= 32'h6A3BCA04;	14'h14F6: data <= 32'h69F1B52D;	14'h14F7: data <= 32'h69A7A057;	14'h14F8: data <= 32'h695D8B80;	14'h14F9: data <= 32'h691376A9;	14'h14FA: data <= 32'h68C961D2;	14'h14FB: data <= 32'h687F4CFB;	14'h14FC: data <= 32'h68353824;	14'h14FD: data <= 32'h67EB234D;	14'h14FE: data <= 32'h67A10E76;	14'h14FF: data <= 32'h6756F99F;	14'h1500: data <= 32'h670CE4C8;	14'h1501: data <= 32'h66C2CFF1;	14'h1502: data <= 32'h6678BB1A;	14'h1503: data <= 32'h662EA643;	14'h1504: data <= 32'h65E4916C;	14'h1505: data <= 32'h659A7C95;	14'h1506: data <= 32'h655067BE;	14'h1507: data <= 32'h650652E7;	14'h1508: data <= 32'h64BC3E11;	14'h1509: data <= 32'h6472293A;	14'h150A: data <= 32'h64281463;	14'h150B: data <= 32'h63DDFF8C;	14'h150C: data <= 32'h6393EAB5;	14'h150D: data <= 32'h6349D5DE;	14'h150E: data <= 32'h62FFC107;	14'h150F: data <= 32'h62B5AC30;	14'h1510: data <= 32'h626B9759;	14'h1511: data <= 32'h62218282;	14'h1512: data <= 32'h61D6E8E5;	14'h1513: data <= 32'h61844545;	14'h1514: data <= 32'h6131A1A5;	14'h1515: data <= 32'h60DEFE05;	14'h1516: data <= 32'h608C5A65;	14'h1517: data <= 32'h6039B6C6;	14'h1518: data <= 32'h5FE71326;	14'h1519: data <= 32'h5F946F86;	14'h151A: data <= 32'h5F41CBE6;	14'h151B: data <= 32'h5EEF2846;	14'h151C: data <= 32'h5E9C84A6;	14'h151D: data <= 32'h5E49E106;	14'h151E: data <= 32'h5DF73D67;	14'h151F: data <= 32'h5DA499C7;	14'h1520: data <= 32'h5D51F627;	14'h1521: data <= 32'h5CFF5287;	14'h1522: data <= 32'h5CACAEE7;	14'h1523: data <= 32'h5C5A0B47;	14'h1524: data <= 32'h5C0767A8;	14'h1525: data <= 32'h5BB4C408;	14'h1526: data <= 32'h5B622068;	14'h1527: data <= 32'h5B0F7CC8;	14'h1528: data <= 32'h5ABCD928;	14'h1529: data <= 32'h5A6A3588;	14'h152A: data <= 32'h5A1791E8;	14'h152B: data <= 32'h59C4EE49;	14'h152C: data <= 32'h59724AA9;	14'h152D: data <= 32'h591FA709;	14'h152E: data <= 32'h58CD0369;	14'h152F: data <= 32'h587A5FC9;	14'h1530: data <= 32'h5827BC29;	14'h1531: data <= 32'h57D1D04C;	14'h1532: data <= 32'h577AD78D;	14'h1533: data <= 32'h5723DECF;	14'h1534: data <= 32'h56CCE610;	14'h1535: data <= 32'h5675ED52;	14'h1536: data <= 32'h561EF494;	14'h1537: data <= 32'h55C7FBD5;	14'h1538: data <= 32'h55710317;	14'h1539: data <= 32'h551A0A58;	14'h153A: data <= 32'h54C3119A;	14'h153B: data <= 32'h546C18DC;	14'h153C: data <= 32'h5415201D;	14'h153D: data <= 32'h53BE275F;	14'h153E: data <= 32'h53672EA1;	14'h153F: data <= 32'h531035E2;	14'h1540: data <= 32'h52B93D24;	14'h1541: data <= 32'h52624465;	14'h1542: data <= 32'h520B4BA7;	14'h1543: data <= 32'h51B452E9;	14'h1544: data <= 32'h515D5A2A;	14'h1545: data <= 32'h5106616C;	14'h1546: data <= 32'h50AF68AD;	14'h1547: data <= 32'h50586FEF;	14'h1548: data <= 32'h50017731;	14'h1549: data <= 32'h4FAA7E72;	14'h154A: data <= 32'h4F5385B4;	14'h154B: data <= 32'h4EFC8CF6;	14'h154C: data <= 32'h4EA59437;	14'h154D: data <= 32'h4E4E9B79;	14'h154E: data <= 32'h4DF7A2BA;	14'h154F: data <= 32'h4DA0A9FC;	14'h1550: data <= 32'h4D49B13E;	14'h1551: data <= 32'h4CF2B87F;	14'h1552: data <= 32'h4C9BBFC1;	14'h1553: data <= 32'h4C44C703;	14'h1554: data <= 32'h4BEDCE44;	14'h1555: data <= 32'h4B96D586;	14'h1556: data <= 32'h4B3FDCC7;	14'h1557: data <= 32'h4AE8E409;	14'h1558: data <= 32'h4A91EB4B;	14'h1559: data <= 32'h4A3AF28C;	14'h155A: data <= 32'h49E3F9CE;	14'h155B: data <= 32'h498D0110;	14'h155C: data <= 32'h49360851;	14'h155D: data <= 32'h48DF0F93;	14'h155E: data <= 32'h488816D5;	14'h155F: data <= 32'h48311E16;	14'h1560: data <= 32'h47DA2558;	14'h1561: data <= 32'h47832C9A;	14'h1562: data <= 32'h472C33DB;	14'h1563: data <= 32'h46D53B1D;	14'h1564: data <= 32'h467E425F;	14'h1565: data <= 32'h462749A0;	14'h1566: data <= 32'h45D050E2;	14'h1567: data <= 32'h45795823;	14'h1568: data <= 32'h45225F65;	14'h1569: data <= 32'h44CB66A7;	14'h156A: data <= 32'h44746DE8;	14'h156B: data <= 32'h441D752A;	14'h156C: data <= 32'h43C67C6C;	14'h156D: data <= 32'h43702293;	14'h156E: data <= 32'h431D428D;	14'h156F: data <= 32'h42CA6288;	14'h1570: data <= 32'h42778282;	14'h1571: data <= 32'h4224A27C;	14'h1572: data <= 32'h41D1C277;	14'h1573: data <= 32'h417EE271;	14'h1574: data <= 32'h412C026C;	14'h1575: data <= 32'h40D92266;	14'h1576: data <= 32'h40864260;	14'h1577: data <= 32'h4033625B;	14'h1578: data <= 32'h3FE08255;	14'h1579: data <= 32'h3F8DA24F;	14'h157A: data <= 32'h3F3AC24A;	14'h157B: data <= 32'h3EE7E244;	14'h157C: data <= 32'h3E95023F;	14'h157D: data <= 32'h3E422239;	14'h157E: data <= 32'h3DEF4233;	14'h157F: data <= 32'h3D9C622E;	14'h1580: data <= 32'h3D498228;	14'h1581: data <= 32'h3CF6A222;	14'h1582: data <= 32'h3CA3C21D;	14'h1583: data <= 32'h3C50E217;	14'h1584: data <= 32'h3BFE0211;	14'h1585: data <= 32'h3BAB220C;	14'h1586: data <= 32'h3B584206;	14'h1587: data <= 32'h3B056201;	14'h1588: data <= 32'h3AB281FB;	14'h1589: data <= 32'h3A5FA1F5;	14'h158A: data <= 32'h3A0CC1F0;	14'h158B: data <= 32'h39B9E1EA;	14'h158C: data <= 32'h396DE2E8;	14'h158D: data <= 32'h39231E5D;	14'h158E: data <= 32'h38D859D3;	14'h158F: data <= 32'h388D9548;	14'h1590: data <= 32'h3842D0BD;	14'h1591: data <= 32'h37F80C33;	14'h1592: data <= 32'h37AD47A8;	14'h1593: data <= 32'h3762831D;	14'h1594: data <= 32'h3717BE93;	14'h1595: data <= 32'h36CCFA08;	14'h1596: data <= 32'h3682357D;	14'h1597: data <= 32'h363770F3;	14'h1598: data <= 32'h35ECAC68;	14'h1599: data <= 32'h35A1E7DD;	14'h159A: data <= 32'h35572353;	14'h159B: data <= 32'h350C5EC8;	14'h159C: data <= 32'h34C19A3D;	14'h159D: data <= 32'h3476D5B3;	14'h159E: data <= 32'h342C1128;	14'h159F: data <= 32'h33E14C9D;	14'h15A0: data <= 32'h33968813;	14'h15A1: data <= 32'h334BC388;	14'h15A2: data <= 32'h3300FEFD;	14'h15A3: data <= 32'h32B63A73;	14'h15A4: data <= 32'h326B75E8;	14'h15A5: data <= 32'h3220B15D;	14'h15A6: data <= 32'h31D5ECD3;	14'h15A7: data <= 32'h318B2848;	14'h15A8: data <= 32'h314063BD;	14'h15A9: data <= 32'h30F59F33;	14'h15AA: data <= 32'h30B116F3;	14'h15AB: data <= 32'h3071C0F2;	14'h15AC: data <= 32'h30326AF1;	14'h15AD: data <= 32'h2FF314F0;	14'h15AE: data <= 32'h2FB3BEEE;	14'h15AF: data <= 32'h2F7468ED;	14'h15B0: data <= 32'h2F3512EC;	14'h15B1: data <= 32'h2EF5BCEB;	14'h15B2: data <= 32'h2EB666EA;	14'h15B3: data <= 32'h2E7710E9;	14'h15B4: data <= 32'h2E37BAE8;	14'h15B5: data <= 32'h2DF864E7;	14'h15B6: data <= 32'h2DB90EE6;	14'h15B7: data <= 32'h2D79B8E4;	14'h15B8: data <= 32'h2D3A62E3;	14'h15B9: data <= 32'h2CFB0CE2;	14'h15BA: data <= 32'h2CBBB6E1;	14'h15BB: data <= 32'h2C7C60E0;	14'h15BC: data <= 32'h2C3D0ADF;	14'h15BD: data <= 32'h2BFDB4DE;	14'h15BE: data <= 32'h2BBE5EDD;	14'h15BF: data <= 32'h2B7F08DC;	14'h15C0: data <= 32'h2B3FB2DA;	14'h15C1: data <= 32'h2B005CD9;	14'h15C2: data <= 32'h2AC106D8;	14'h15C3: data <= 32'h2A81B0D7;	14'h15C4: data <= 32'h2A425AD6;	14'h15C5: data <= 32'h2A0304D5;	14'h15C6: data <= 32'h29C3AED4;	14'h15C7: data <= 32'h298458D3;	14'h15C8: data <= 32'h2948500D;	14'h15C9: data <= 32'h291698A3;	14'h15CA: data <= 32'h28E4E138;	14'h15CB: data <= 32'h28B329CD;	14'h15CC: data <= 32'h28817262;	14'h15CD: data <= 32'h284FBAF7;	14'h15CE: data <= 32'h281E038D;	14'h15CF: data <= 32'h27EC4C22;	14'h15D0: data <= 32'h27BA94B7;	14'h15D1: data <= 32'h2788DD4C;	14'h15D2: data <= 32'h275725E2;	14'h15D3: data <= 32'h27256E77;	14'h15D4: data <= 32'h26F3B70C;	14'h15D5: data <= 32'h26C1FFA1;	14'h15D6: data <= 32'h26904837;	14'h15D7: data <= 32'h265E90CC;	14'h15D8: data <= 32'h262CD961;	14'h15D9: data <= 32'h25FB21F6;	14'h15DA: data <= 32'h25C96A8B;	14'h15DB: data <= 32'h2597B321;	14'h15DC: data <= 32'h2565FBB6;	14'h15DD: data <= 32'h2534444B;	14'h15DE: data <= 32'h25028CE0;	14'h15DF: data <= 32'h24D0D576;	14'h15E0: data <= 32'h249F1E0B;	14'h15E1: data <= 32'h246D66A0;	14'h15E2: data <= 32'h243BAF35;	14'h15E3: data <= 32'h2409F7CB;	14'h15E4: data <= 32'h23D84060;	14'h15E5: data <= 32'h23A688F5;	14'h15E6: data <= 32'h2374D18A;	14'h15E7: data <= 32'h23512F82;	14'h15E8: data <= 32'h232E7616;	14'h15E9: data <= 32'h230BBCA9;	14'h15EA: data <= 32'h22E9033C;	14'h15EB: data <= 32'h22C649CF;	14'h15EC: data <= 32'h22A39062;	14'h15ED: data <= 32'h2280D6F5;	14'h15EE: data <= 32'h225E1D88;	14'h15EF: data <= 32'h223B641B;	14'h15F0: data <= 32'h2218AAAF;	14'h15F1: data <= 32'h21F5F142;	14'h15F2: data <= 32'h21D337D5;	14'h15F3: data <= 32'h21B07E68;	14'h15F4: data <= 32'h218DC4FB;	14'h15F5: data <= 32'h216B0B8E;	14'h15F6: data <= 32'h21485221;	14'h15F7: data <= 32'h212598B4;	14'h15F8: data <= 32'h2102DF48;	14'h15F9: data <= 32'h20E025DB;	14'h15FA: data <= 32'h20BD6C6E;	14'h15FB: data <= 32'h209AB301;	14'h15FC: data <= 32'h2077F994;	14'h15FD: data <= 32'h20554027;	14'h15FE: data <= 32'h203286BA;	14'h15FF: data <= 32'h200FCD4E;	14'h1600: data <= 32'h1FED13E1;	14'h1601: data <= 32'h1FCA5A74;	14'h1602: data <= 32'h1FA7A107;	14'h1603: data <= 32'h1F84E79A;	14'h1604: data <= 32'h1F622E2D;	14'h1605: data <= 32'h1F48E6A7;	14'h1606: data <= 32'h1F3504C8;	14'h1607: data <= 32'h1F2122EA;	14'h1608: data <= 32'h1F0D410B;	14'h1609: data <= 32'h1EF95F2D;	14'h160A: data <= 32'h1EE57D4F;	14'h160B: data <= 32'h1ED19B70;	14'h160C: data <= 32'h1EBDB992;	14'h160D: data <= 32'h1EA9D7B4;	14'h160E: data <= 32'h1E95F5D5;	14'h160F: data <= 32'h1E8213F7;	14'h1610: data <= 32'h1E6E3218;	14'h1611: data <= 32'h1E5A503A;	14'h1612: data <= 32'h1E466E5C;	14'h1613: data <= 32'h1E328C7D;	14'h1614: data <= 32'h1E1EAA9F;	14'h1615: data <= 32'h1E0AC8C0;	14'h1616: data <= 32'h1DF6E6E2;	14'h1617: data <= 32'h1DE30504;	14'h1618: data <= 32'h1DCF2325;	14'h1619: data <= 32'h1DBB4147;	14'h161A: data <= 32'h1DA75F69;	14'h161B: data <= 32'h1D937D8A;	14'h161C: data <= 32'h1D7F9BAC;	14'h161D: data <= 32'h1D6BB9CD;	14'h161E: data <= 32'h1D57D7EF;	14'h161F: data <= 32'h1D43F611;	14'h1620: data <= 32'h1D301432;	14'h1621: data <= 32'h1D1C3254;	14'h1622: data <= 32'h1D085075;	14'h1623: data <= 32'h1CF88EA2;	14'h1624: data <= 32'h1CF10CE4;	14'h1625: data <= 32'h1CE98B26;	14'h1626: data <= 32'h1CE20969;	14'h1627: data <= 32'h1CDA87AB;	14'h1628: data <= 32'h1CD305ED;	14'h1629: data <= 32'h1CCB8430;	14'h162A: data <= 32'h1CC40272;	14'h162B: data <= 32'h1CBC80B4;	14'h162C: data <= 32'h1CB4FEF6;	14'h162D: data <= 32'h1CAD7D39;	14'h162E: data <= 32'h1CA5FB7B;	14'h162F: data <= 32'h1C9E79BD;	14'h1630: data <= 32'h1C96F800;	14'h1631: data <= 32'h1C8F7642;	14'h1632: data <= 32'h1C87F484;	14'h1633: data <= 32'h1C8072C6;	14'h1634: data <= 32'h1C78F109;	14'h1635: data <= 32'h1C716F4B;	14'h1636: data <= 32'h1C69ED8D;	14'h1637: data <= 32'h1C626BD0;	14'h1638: data <= 32'h1C5AEA12;	14'h1639: data <= 32'h1C536854;	14'h163A: data <= 32'h1C4BE696;	14'h163B: data <= 32'h1C4464D9;	14'h163C: data <= 32'h1C3CE31B;	14'h163D: data <= 32'h1C35615D;	14'h163E: data <= 32'h1C2DDFA0;	14'h163F: data <= 32'h1C265DE2;	14'h1640: data <= 32'h1C1EDC24;	14'h1641: data <= 32'h1C1799A0;	14'h1642: data <= 32'h1C183E59;	14'h1643: data <= 32'h1C18E311;	14'h1644: data <= 32'h1C1987CA;	14'h1645: data <= 32'h1C1A2C82;	14'h1646: data <= 32'h1C1AD13B;	14'h1647: data <= 32'h1C1B75F3;	14'h1648: data <= 32'h1C1C1AAC;	14'h1649: data <= 32'h1C1CBF64;	14'h164A: data <= 32'h1C1D641D;	14'h164B: data <= 32'h1C1E08D5;	14'h164C: data <= 32'h1C1EAD8E;	14'h164D: data <= 32'h1C1F5246;	14'h164E: data <= 32'h1C1FF6FF;	14'h164F: data <= 32'h1C209BB7;	14'h1650: data <= 32'h1C214070;	14'h1651: data <= 32'h1C21E528;	14'h1652: data <= 32'h1C2289E1;	14'h1653: data <= 32'h1C232E99;	14'h1654: data <= 32'h1C23D352;	14'h1655: data <= 32'h1C24780A;	14'h1656: data <= 32'h1C251CC3;	14'h1657: data <= 32'h1C25C17B;	14'h1658: data <= 32'h1C266634;	14'h1659: data <= 32'h1C270AEC;	14'h165A: data <= 32'h1C27AFA5;	14'h165B: data <= 32'h1C28545D;	14'h165C: data <= 32'h1C28F916;	14'h165D: data <= 32'h1C299DCE;	14'h165E: data <= 32'h1C2A4287;	14'h165F: data <= 32'h1C2AE73F;	14'h1660: data <= 32'h1C2E2ED3;	14'h1661: data <= 32'h1C327378;	14'h1662: data <= 32'h1C36B81E;	14'h1663: data <= 32'h1C3AFCC3;	14'h1664: data <= 32'h1C3F4169;	14'h1665: data <= 32'h1C43860F;	14'h1666: data <= 32'h1C47CAB4;	14'h1667: data <= 32'h1C4C0F5A;	14'h1668: data <= 32'h1C505400;	14'h1669: data <= 32'h1C5498A5;	14'h166A: data <= 32'h1C58DD4B;	14'h166B: data <= 32'h1C5D21F1;	14'h166C: data <= 32'h1C616696;	14'h166D: data <= 32'h1C65AB3C;	14'h166E: data <= 32'h1C69EFE1;	14'h166F: data <= 32'h1C6E3487;	14'h1670: data <= 32'h1C72792D;	14'h1671: data <= 32'h1C76BDD2;	14'h1672: data <= 32'h1C7B0278;	14'h1673: data <= 32'h1C7F471E;	14'h1674: data <= 32'h1C838BC3;	14'h1675: data <= 32'h1C87D069;	14'h1676: data <= 32'h1C8C150F;	14'h1677: data <= 32'h1C9059B4;	14'h1678: data <= 32'h1C949E5A;	14'h1679: data <= 32'h1C98E2FF;	14'h167A: data <= 32'h1C9D27A5;	14'h167B: data <= 32'h1CA16C4B;	14'h167C: data <= 32'h1CA5B0F0;	14'h167D: data <= 32'h1CA9F596;	14'h167E: data <= 32'h1CADBA1E;	14'h167F: data <= 32'h1CB0D0C7;	14'h1680: data <= 32'h1CB3E76F;	14'h1681: data <= 32'h1CB6FE18;	14'h1682: data <= 32'h1CBA14C1;	14'h1683: data <= 32'h1CBD2B6A;	14'h1684: data <= 32'h1CC04212;	14'h1685: data <= 32'h1CC358BB;	14'h1686: data <= 32'h1CC66F64;	14'h1687: data <= 32'h1CC9860D;	14'h1688: data <= 32'h1CCC9CB6;	14'h1689: data <= 32'h1CCFB35E;	14'h168A: data <= 32'h1CD2CA07;	14'h168B: data <= 32'h1CD5E0B0;	14'h168C: data <= 32'h1CD8F759;	14'h168D: data <= 32'h1CDC0E01;	14'h168E: data <= 32'h1CDF24AA;	14'h168F: data <= 32'h1CE23B53;	14'h1690: data <= 32'h1CE551FC;	14'h1691: data <= 32'h1CE868A4;	14'h1692: data <= 32'h1CEB7F4D;	14'h1693: data <= 32'h1CEE95F6;	14'h1694: data <= 32'h1CF1AC9F;	14'h1695: data <= 32'h1CF4C348;	14'h1696: data <= 32'h1CF7D9F0;	14'h1697: data <= 32'h1CFAF099;	14'h1698: data <= 32'h1CFE0742;	14'h1699: data <= 32'h1D011DEB;	14'h169A: data <= 32'h1D043493;	14'h169B: data <= 32'h1D074B3C;	14'h169C: data <= 32'h1D09A437;	14'h169D: data <= 32'h1D069E07;	14'h169E: data <= 32'h1D0397D7;	14'h169F: data <= 32'h1D0091A8;	14'h16A0: data <= 32'h1CFD8B78;	14'h16A1: data <= 32'h1CFA8548;	14'h16A2: data <= 32'h1CF77F18;	14'h16A3: data <= 32'h1CF478E8;	14'h16A4: data <= 32'h1CF172B8;	14'h16A5: data <= 32'h1CEE6C88;	14'h16A6: data <= 32'h1CEB6658;	14'h16A7: data <= 32'h1CE86028;	14'h16A8: data <= 32'h1CE559F9;	14'h16A9: data <= 32'h1CE253C9;	14'h16AA: data <= 32'h1CDF4D99;	14'h16AB: data <= 32'h1CDC4769;	14'h16AC: data <= 32'h1CD94139;	14'h16AD: data <= 32'h1CD63B09;	14'h16AE: data <= 32'h1CD334D9;	14'h16AF: data <= 32'h1CD02EA9;	14'h16B0: data <= 32'h1CCD2879;	14'h16B1: data <= 32'h1CCA2249;	14'h16B2: data <= 32'h1CC71C1A;	14'h16B3: data <= 32'h1CC415EA;	14'h16B4: data <= 32'h1CC10FBA;	14'h16B5: data <= 32'h1CBE098A;	14'h16B6: data <= 32'h1CBB035A;	14'h16B7: data <= 32'h1CB7FD2A;	14'h16B8: data <= 32'h1CB4F6FA;	14'h16B9: data <= 32'h1CB1F0CA;	14'h16BA: data <= 32'h1CAEEA9A;	14'h16BB: data <= 32'h1CA407D4;	14'h16BC: data <= 32'h1C9765D0;	14'h16BD: data <= 32'h1C8AC3CC;	14'h16BE: data <= 32'h1C7E21C8;	14'h16BF: data <= 32'h1C717FC4;	14'h16C0: data <= 32'h1C64DDC0;	14'h16C1: data <= 32'h1C583BBC;	14'h16C2: data <= 32'h1C4B99B8;	14'h16C3: data <= 32'h1C3EF7B4;	14'h16C4: data <= 32'h1C3255B0;	14'h16C5: data <= 32'h1C25B3AC;	14'h16C6: data <= 32'h1C1911A8;	14'h16C7: data <= 32'h1C0C6FA3;	14'h16C8: data <= 32'h1BFFCD9F;	14'h16C9: data <= 32'h1BF32B9B;	14'h16CA: data <= 32'h1BE68997;	14'h16CB: data <= 32'h1BD9E793;	14'h16CC: data <= 32'h1BCD458F;	14'h16CD: data <= 32'h1BC0A38B;	14'h16CE: data <= 32'h1BB40187;	14'h16CF: data <= 32'h1BA75F83;	14'h16D0: data <= 32'h1B9ABD7F;	14'h16D1: data <= 32'h1B8E1B7B;	14'h16D2: data <= 32'h1B817977;	14'h16D3: data <= 32'h1B74D773;	14'h16D4: data <= 32'h1B68356F;	14'h16D5: data <= 32'h1B5B936B;	14'h16D6: data <= 32'h1B4EF167;	14'h16D7: data <= 32'h1B424F63;	14'h16D8: data <= 32'h1B35AD5E;	14'h16D9: data <= 32'h1B235500;	14'h16DA: data <= 32'h1B0B9C4C;	14'h16DB: data <= 32'h1AF3E399;	14'h16DC: data <= 32'h1ADC2AE5;	14'h16DD: data <= 32'h1AC47231;	14'h16DE: data <= 32'h1AACB97E;	14'h16DF: data <= 32'h1A9500CA;	14'h16E0: data <= 32'h1A7D4816;	14'h16E1: data <= 32'h1A658F62;	14'h16E2: data <= 32'h1A4DD6AF;	14'h16E3: data <= 32'h1A361DFB;	14'h16E4: data <= 32'h1A1E6547;	14'h16E5: data <= 32'h1A06AC94;	14'h16E6: data <= 32'h19EEF3E0;	14'h16E7: data <= 32'h19D73B2C;	14'h16E8: data <= 32'h19BF8279;	14'h16E9: data <= 32'h19A7C9C5;	14'h16EA: data <= 32'h19901111;	14'h16EB: data <= 32'h1978585E;	14'h16EC: data <= 32'h19609FAA;	14'h16ED: data <= 32'h1948E6F6;	14'h16EE: data <= 32'h19312E43;	14'h16EF: data <= 32'h1919758F;	14'h16F0: data <= 32'h1901BCDB;	14'h16F1: data <= 32'h18EA0427;	14'h16F2: data <= 32'h18D24B74;	14'h16F3: data <= 32'h18BA92C0;	14'h16F4: data <= 32'h18A2DA0C;	14'h16F5: data <= 32'h188B2159;	14'h16F6: data <= 32'h187368A5;	14'h16F7: data <= 32'h1859432A;	14'h16F8: data <= 32'h18361BEC;	14'h16F9: data <= 32'h1812F4AF;	14'h16FA: data <= 32'h17EFCD72;	14'h16FB: data <= 32'h17CCA635;	14'h16FC: data <= 32'h17A97EF7;	14'h16FD: data <= 32'h178657BA;	14'h16FE: data <= 32'h1763307D;	14'h16FF: data <= 32'h17400940;	14'h1700: data <= 32'h171CE202;	14'h1701: data <= 32'h16F9BAC5;	14'h1702: data <= 32'h16D69388;	14'h1703: data <= 32'h16B36C4B;	14'h1704: data <= 32'h1690450D;	14'h1705: data <= 32'h166D1DD0;	14'h1706: data <= 32'h1649F693;	14'h1707: data <= 32'h1626CF56;	14'h1708: data <= 32'h1603A818;	14'h1709: data <= 32'h15E080DB;	14'h170A: data <= 32'h15BD599E;	14'h170B: data <= 32'h159A3261;	14'h170C: data <= 32'h15770B23;	14'h170D: data <= 32'h1553E3E6;	14'h170E: data <= 32'h1530BCA9;	14'h170F: data <= 32'h150D956C;	14'h1710: data <= 32'h14EA6E2F;	14'h1711: data <= 32'h14C746F1;	14'h1712: data <= 32'h14A41FB4;	14'h1713: data <= 32'h1480F877;	14'h1714: data <= 32'h145DD13A;	14'h1715: data <= 32'h143AA9FC;	14'h1716: data <= 32'h140DEAE9;	14'h1717: data <= 32'h13E03641;	14'h1718: data <= 32'h13B28198;	14'h1719: data <= 32'h1384CCF0;	14'h171A: data <= 32'h13571847;	14'h171B: data <= 32'h1329639F;	14'h171C: data <= 32'h12FBAEF6;	14'h171D: data <= 32'h12CDFA4E;	14'h171E: data <= 32'h12A045A5;	14'h171F: data <= 32'h127290FD;	14'h1720: data <= 32'h1244DC54;	14'h1721: data <= 32'h121727AC;	14'h1722: data <= 32'h11E97303;	14'h1723: data <= 32'h11BBBE5B;	14'h1724: data <= 32'h118E09B2;	14'h1725: data <= 32'h1160550A;	14'h1726: data <= 32'h1132A061;	14'h1727: data <= 32'h1104EBB9;	14'h1728: data <= 32'h10D73710;	14'h1729: data <= 32'h10A98268;	14'h172A: data <= 32'h107BCDC0;	14'h172B: data <= 32'h104E1917;	14'h172C: data <= 32'h1020646F;	14'h172D: data <= 32'h0FF2AFC6;	14'h172E: data <= 32'h0FC4FB1E;	14'h172F: data <= 32'h0F974675;	14'h1730: data <= 32'h0F6991CD;	14'h1731: data <= 32'h0F3BDD24;	14'h1732: data <= 32'h0F0E287C;	14'h1733: data <= 32'h0EE073D3;	14'h1734: data <= 32'h0EAE0A8B;	14'h1735: data <= 32'h0E789241;	14'h1736: data <= 32'h0E4319F8;	14'h1737: data <= 32'h0E0DA1AE;	14'h1738: data <= 32'h0DD82965;	14'h1739: data <= 32'h0DA2B11B;	14'h173A: data <= 32'h0D6D38D1;	14'h173B: data <= 32'h0D37C088;	14'h173C: data <= 32'h0D02483E;	14'h173D: data <= 32'h0CCCCFF5;	14'h173E: data <= 32'h0C9757AB;	14'h173F: data <= 32'h0C61DF61;	14'h1740: data <= 32'h0C2C6718;	14'h1741: data <= 32'h0BF6EECE;	14'h1742: data <= 32'h0BC17685;	14'h1743: data <= 32'h0B8BFE3B;	14'h1744: data <= 32'h0B5685F2;	14'h1745: data <= 32'h0B210DA8;	14'h1746: data <= 32'h0AEB955E;	14'h1747: data <= 32'h0AB61D15;	14'h1748: data <= 32'h0A80A4CB;	14'h1749: data <= 32'h0A4B2C82;	14'h174A: data <= 32'h0A15B438;	14'h174B: data <= 32'h09E03BEE;	14'h174C: data <= 32'h09AAC3A5;	14'h174D: data <= 32'h09754B5B;	14'h174E: data <= 32'h093FD312;	14'h174F: data <= 32'h090A5AC8;	14'h1750: data <= 32'h08D4E27E;	14'h1751: data <= 32'h089F6A35;	14'h1752: data <= 32'h0865CFB7;	14'h1753: data <= 32'h0822B359;	14'h1754: data <= 32'h07DF96FB;	14'h1755: data <= 32'h079C7A9E;	14'h1756: data <= 32'h07595E40;	14'h1757: data <= 32'h071641E3;	14'h1758: data <= 32'h06D32585;	14'h1759: data <= 32'h06900927;	14'h175A: data <= 32'h064CECCA;	14'h175B: data <= 32'h0609D06C;	14'h175C: data <= 32'h05C6B40F;	14'h175D: data <= 32'h058397B1;	14'h175E: data <= 32'h05407B53;	14'h175F: data <= 32'h04FD5EF6;	14'h1760: data <= 32'h04BA4298;	14'h1761: data <= 32'h0477263B;	14'h1762: data <= 32'h043409DD;	14'h1763: data <= 32'h03F0ED7F;	14'h1764: data <= 32'h03ADD122;	14'h1765: data <= 32'h036AB4C4;	14'h1766: data <= 32'h03279867;	14'h1767: data <= 32'h02E47C09;	14'h1768: data <= 32'h02A15FAB;	14'h1769: data <= 32'h025E434E;	14'h176A: data <= 32'h021B26F0;	14'h176B: data <= 32'h01D80A93;	14'h176C: data <= 32'h0194EE35;	14'h176D: data <= 32'h0151D1D7;	14'h176E: data <= 32'h010EB57A;	14'h176F: data <= 32'h00CB991C;	14'h1770: data <= 32'hE67EEA69;	14'h1771: data <= 32'hE6993A35;	14'h1772: data <= 32'hE6B38A00;	14'h1773: data <= 32'hE6CDD9CB;	14'h1774: data <= 32'hE6E82996;	14'h1775: data <= 32'hE7027961;	14'h1776: data <= 32'hE71CC92D;	14'h1777: data <= 32'hE73718F8;	14'h1778: data <= 32'hE75168C3;	14'h1779: data <= 32'hE76BB88E;	14'h177A: data <= 32'hE7860859;	14'h177B: data <= 32'hE7A05824;	14'h177C: data <= 32'hE7BAA7F0;	14'h177D: data <= 32'hE7D4F7BB;	14'h177E: data <= 32'hE7EF4786;	14'h177F: data <= 32'hE8099751;	14'h1780: data <= 32'hE823E71C;	14'h1781: data <= 32'hE83E36E8;	14'h1782: data <= 32'hE85886B3;	14'h1783: data <= 32'hE872D67E;	14'h1784: data <= 32'hE88D2649;	14'h1785: data <= 32'hE8A77614;	14'h1786: data <= 32'hE8C1C5DF;	14'h1787: data <= 32'hE8DC15AB;	14'h1788: data <= 32'hE8F66576;	14'h1789: data <= 32'hE910B541;	14'h178A: data <= 32'hE92B050C;	14'h178B: data <= 32'hE94554D7;	14'h178C: data <= 32'hE95FA4A3;	14'h178D: data <= 32'hE979F46E;	14'h178E: data <= 32'hE9944439;	14'h178F: data <= 32'hE9AE9404;	14'h1790: data <= 32'hE9C8E3CF;	14'h1791: data <= 32'hE9E3339A;	14'h1792: data <= 32'hE9FD8366;	14'h1793: data <= 32'hEA17D331;	14'h1794: data <= 32'hEA3222FC;	14'h1795: data <= 32'hEA495186;	14'h1796: data <= 32'hEA5FF8A3;	14'h1797: data <= 32'hEA769FC0;	14'h1798: data <= 32'hEA8D46DD;	14'h1799: data <= 32'hEAA3EDFB;	14'h179A: data <= 32'hEABA9518;	14'h179B: data <= 32'hEAD13C35;	14'h179C: data <= 32'hEAE7E353;	14'h179D: data <= 32'hEAFE8A70;	14'h179E: data <= 32'hEB15318D;	14'h179F: data <= 32'hEB2BD8AA;	14'h17A0: data <= 32'hEB427FC8;	14'h17A1: data <= 32'hEB5926E5;	14'h17A2: data <= 32'hEB6FCE02;	14'h17A3: data <= 32'hEB867520;	14'h17A4: data <= 32'hEB9D1C3D;	14'h17A5: data <= 32'hEBB3C35A;	14'h17A6: data <= 32'hEBCA6A77;	14'h17A7: data <= 32'hEBE11195;	14'h17A8: data <= 32'hEBF7B8B2;	14'h17A9: data <= 32'hEC0E5FCF;	14'h17AA: data <= 32'hEC2506EC;	14'h17AB: data <= 32'hEC3BAE0A;	14'h17AC: data <= 32'hEC525527;	14'h17AD: data <= 32'hEC68FC44;	14'h17AE: data <= 32'hEC7FA362;	14'h17AF: data <= 32'hEC964A7F;	14'h17B0: data <= 32'hECACF19C;	14'h17B1: data <= 32'hECC398B9;	14'h17B2: data <= 32'hECDA3FD7;	14'h17B3: data <= 32'hECF0E6F4;	14'h17B4: data <= 32'hED078E11;	14'h17B5: data <= 32'hED1E352E;	14'h17B6: data <= 32'hED34DC4C;	14'h17B7: data <= 32'hED4B8369;	14'h17B8: data <= 32'hED622A86;	14'h17B9: data <= 32'hED7649A1;	14'h17BA: data <= 32'hED896122;	14'h17BB: data <= 32'hED9C78A3;	14'h17BC: data <= 32'hEDAF9024;	14'h17BD: data <= 32'hEDC2A7A6;	14'h17BE: data <= 32'hEDD5BF27;	14'h17BF: data <= 32'hEDE8D6A8;	14'h17C0: data <= 32'hEDFBEE29;	14'h17C1: data <= 32'hEE0F05AB;	14'h17C2: data <= 32'hEE221D2C;	14'h17C3: data <= 32'hEE3534AD;	14'h17C4: data <= 32'hEE484C2F;	14'h17C5: data <= 32'hEE5B63B0;	14'h17C6: data <= 32'hEE6E7B31;	14'h17C7: data <= 32'hEE8192B2;	14'h17C8: data <= 32'hEE94AA34;	14'h17C9: data <= 32'hEEA7C1B5;	14'h17CA: data <= 32'hEEBAD936;	14'h17CB: data <= 32'hEECDF0B7;	14'h17CC: data <= 32'hEEE10839;	14'h17CD: data <= 32'hEEF41FBA;	14'h17CE: data <= 32'hEF07373B;	14'h17CF: data <= 32'hEF1A4EBC;	14'h17D0: data <= 32'hEF2D663E;	14'h17D1: data <= 32'hEF407DBF;	14'h17D2: data <= 32'hEF539540;	14'h17D3: data <= 32'hEF66ACC1;	14'h17D4: data <= 32'hEF79C443;	14'h17D5: data <= 32'hEF8CDBC4;	14'h17D6: data <= 32'hEF9FF345;	14'h17D7: data <= 32'hEFB30AC6;	14'h17D8: data <= 32'hEFC62248;	14'h17D9: data <= 32'hEFD939C9;	14'h17DA: data <= 32'hEFEC514A;	14'h17DB: data <= 32'hEFFF68CC;	14'h17DC: data <= 32'hF012804D;	14'h17DD: data <= 32'hF0242310;	14'h17DE: data <= 32'hF034A851;	14'h17DF: data <= 32'hF0452D93;	14'h17E0: data <= 32'hF055B2D4;	14'h17E1: data <= 32'hF0663816;	14'h17E2: data <= 32'hF076BD57;	14'h17E3: data <= 32'hF0874299;	14'h17E4: data <= 32'hF097C7DA;	14'h17E5: data <= 32'hF0A84D1C;	14'h17E6: data <= 32'hF0B8D25D;	14'h17E7: data <= 32'hF0C9579F;	14'h17E8: data <= 32'hF0D9DCE0;	14'h17E9: data <= 32'hF0EA6222;	14'h17EA: data <= 32'hF0FAE763;	14'h17EB: data <= 32'hF10B6CA5;	14'h17EC: data <= 32'hF11BF1E6;	14'h17ED: data <= 32'hF12C7728;	14'h17EE: data <= 32'hF13CFC69;	14'h17EF: data <= 32'hF14D81AB;	14'h17F0: data <= 32'hF15E06EC;	14'h17F1: data <= 32'hF16E8C2D;	14'h17F2: data <= 32'hF17F116F;	14'h17F3: data <= 32'hF18F96B0;	14'h17F4: data <= 32'hF1A01BF2;	14'h17F5: data <= 32'hF1B0A133;	14'h17F6: data <= 32'hF1C12675;	14'h17F7: data <= 32'hF1D1ABB6;	14'h17F8: data <= 32'hF1E230F8;	14'h17F9: data <= 32'hF1F2B639;	14'h17FA: data <= 32'hF2033B7B;	14'h17FB: data <= 32'hF213C0BC;	14'h17FC: data <= 32'hF22445FE;	14'h17FD: data <= 32'hF234CB3F;	14'h17FE: data <= 32'hF2455081;	14'h17FF: data <= 32'hF255D5C2;	14'h1800: data <= 32'hF2665B04;	14'h1801: data <= 32'hF273E12D;	14'h1802: data <= 32'hF27D4B51;	14'h1803: data <= 32'hF286B575;	14'h1804: data <= 32'hF2901F99;	14'h1805: data <= 32'hF29989BD;	14'h1806: data <= 32'hF2A2F3E1;	14'h1807: data <= 32'hF2AC5E05;	14'h1808: data <= 32'hF2B5C82A;	14'h1809: data <= 32'hF2BF324E;	14'h180A: data <= 32'hF2C89C72;	14'h180B: data <= 32'hF2D20696;	14'h180C: data <= 32'hF2DB70BA;	14'h180D: data <= 32'hF2E4DADE;	14'h180E: data <= 32'hF2EE4502;	14'h180F: data <= 32'hF2F7AF26;	14'h1810: data <= 32'hF301194B;	14'h1811: data <= 32'hF30A836F;	14'h1812: data <= 32'hF313ED93;	14'h1813: data <= 32'hF31D57B7;	14'h1814: data <= 32'hF326C1DB;	14'h1815: data <= 32'hF3302BFF;	14'h1816: data <= 32'hF3399623;	14'h1817: data <= 32'hF3430047;	14'h1818: data <= 32'hF34C6A6C;	14'h1819: data <= 32'hF355D490;	14'h181A: data <= 32'hF35F3EB4;	14'h181B: data <= 32'hF368A8D8;	14'h181C: data <= 32'hF37212FC;	14'h181D: data <= 32'hF37B7D20;	14'h181E: data <= 32'hF384E744;	14'h181F: data <= 32'hF38E5169;	14'h1820: data <= 32'hF397BB8D;	14'h1821: data <= 32'hF3A125B1;	14'h1822: data <= 32'hF3AA8FD5;	14'h1823: data <= 32'hF3B3F9F9;	14'h1824: data <= 32'hF3BD641D;	14'h1825: data <= 32'hF3C52E5F;	14'h1826: data <= 32'hF3C8BBB4;	14'h1827: data <= 32'hF3CC490A;	14'h1828: data <= 32'hF3CFD660;	14'h1829: data <= 32'hF3D363B6;	14'h182A: data <= 32'hF3D6F10C;	14'h182B: data <= 32'hF3DA7E62;	14'h182C: data <= 32'hF3DE0BB8;	14'h182D: data <= 32'hF3E1990E;	14'h182E: data <= 32'hF3E52663;	14'h182F: data <= 32'hF3E8B3B9;	14'h1830: data <= 32'hF3EC410F;	14'h1831: data <= 32'hF3EFCE65;	14'h1832: data <= 32'hF3F35BBB;	14'h1833: data <= 32'hF3F6E911;	14'h1834: data <= 32'hF3FA7667;	14'h1835: data <= 32'hF3FE03BD;	14'h1836: data <= 32'hF4019112;	14'h1837: data <= 32'hF4051E68;	14'h1838: data <= 32'hF408ABBE;	14'h1839: data <= 32'hF40C3914;	14'h183A: data <= 32'hF40FC66A;	14'h183B: data <= 32'hF41353C0;	14'h183C: data <= 32'hF416E116;	14'h183D: data <= 32'hF41A6E6C;	14'h183E: data <= 32'hF41DFBC2;	14'h183F: data <= 32'hF4218917;	14'h1840: data <= 32'hF425166D;	14'h1841: data <= 32'hF428A3C3;	14'h1842: data <= 32'hF42C3119;	14'h1843: data <= 32'hF42FBE6F;	14'h1844: data <= 32'hF4334BC5;	14'h1845: data <= 32'hF436D91B;	14'h1846: data <= 32'hF43A6671;	14'h1847: data <= 32'hF43DF3C6;	14'h1848: data <= 32'hF441811C;	14'h1849: data <= 32'hF444B997;	14'h184A: data <= 32'hF445C6A6;	14'h184B: data <= 32'hF446D3B4;	14'h184C: data <= 32'hF447E0C3;	14'h184D: data <= 32'hF448EDD1;	14'h184E: data <= 32'hF449FAE0;	14'h184F: data <= 32'hF44B07EE;	14'h1850: data <= 32'hF44C14FD;	14'h1851: data <= 32'hF44D220B;	14'h1852: data <= 32'hF44E2F1A;	14'h1853: data <= 32'hF44F3C28;	14'h1854: data <= 32'hF4504937;	14'h1855: data <= 32'hF4515646;	14'h1856: data <= 32'hF4526354;	14'h1857: data <= 32'hF4537063;	14'h1858: data <= 32'hF4547D71;	14'h1859: data <= 32'hF4558A80;	14'h185A: data <= 32'hF456978E;	14'h185B: data <= 32'hF457A49D;	14'h185C: data <= 32'hF458B1AB;	14'h185D: data <= 32'hF459BEBA;	14'h185E: data <= 32'hF45ACBC8;	14'h185F: data <= 32'hF45BD8D7;	14'h1860: data <= 32'hF45CE5E6;	14'h1861: data <= 32'hF45DF2F4;	14'h1862: data <= 32'hF45F0003;	14'h1863: data <= 32'hF4600D11;	14'h1864: data <= 32'hF4611A20;	14'h1865: data <= 32'hF462272E;	14'h1866: data <= 32'hF463343D;	14'h1867: data <= 32'hF464414B;	14'h1868: data <= 32'hF4654E5A;	14'h1869: data <= 32'hF4665B68;	14'h186A: data <= 32'hF4676877;	14'h186B: data <= 32'hF4687586;	14'h186C: data <= 32'hF4698294;	14'h186D: data <= 32'hF46A8FA3;	14'h186E: data <= 32'hF46E4AAF;	14'h186F: data <= 32'hF4720E18;	14'h1870: data <= 32'hF475D182;	14'h1871: data <= 32'hF47994EC;	14'h1872: data <= 32'hF47D5856;	14'h1873: data <= 32'hF4811BBF;	14'h1874: data <= 32'hF484DF29;	14'h1875: data <= 32'hF488A293;	14'h1876: data <= 32'hF48C65FD;	14'h1877: data <= 32'hF4902966;	14'h1878: data <= 32'hF493ECD0;	14'h1879: data <= 32'hF497B03A;	14'h187A: data <= 32'hF49B73A3;	14'h187B: data <= 32'hF49F370D;	14'h187C: data <= 32'hF4A2FA77;	14'h187D: data <= 32'hF4A6BDE1;	14'h187E: data <= 32'hF4AA814A;	14'h187F: data <= 32'hF4AE44B4;	14'h1880: data <= 32'hF4B2081E;	14'h1881: data <= 32'hF4B5CB88;	14'h1882: data <= 32'hF4B98EF1;	14'h1883: data <= 32'hF4BD525B;	14'h1884: data <= 32'hF4C115C5;	14'h1885: data <= 32'hF4C4D92E;	14'h1886: data <= 32'hF4C89C98;	14'h1887: data <= 32'hF4CC6002;	14'h1888: data <= 32'hF4D0236C;	14'h1889: data <= 32'hF4D3E6D5;	14'h188A: data <= 32'hF4D7AA3F;	14'h188B: data <= 32'hF4DB6DA9;	14'h188C: data <= 32'hF4DF3112;	14'h188D: data <= 32'hF4E2F47C;	14'h188E: data <= 32'hF4E6B7E6;	14'h188F: data <= 32'hF4EA7B50;	14'h1890: data <= 32'hF4EE3EB9;	14'h1891: data <= 32'hF4F20223;	14'h1892: data <= 32'hF4F7B66A;	14'h1893: data <= 32'hF4FDC6F8;	14'h1894: data <= 32'hF503D786;	14'h1895: data <= 32'hF509E814;	14'h1896: data <= 32'hF50FF8A2;	14'h1897: data <= 32'hF516092F;	14'h1898: data <= 32'hF51C19BD;	14'h1899: data <= 32'hF5222A4B;	14'h189A: data <= 32'hF5283AD9;	14'h189B: data <= 32'hF52E4B66;	14'h189C: data <= 32'hF5345BF4;	14'h189D: data <= 32'hF53A6C82;	14'h189E: data <= 32'hF5407D10;	14'h189F: data <= 32'hF5468D9E;	14'h18A0: data <= 32'hF54C9E2B;	14'h18A1: data <= 32'hF552AEB9;	14'h18A2: data <= 32'hF558BF47;	14'h18A3: data <= 32'hF55ECFD5;	14'h18A4: data <= 32'hF564E062;	14'h18A5: data <= 32'hF56AF0F0;	14'h18A6: data <= 32'hF571017E;	14'h18A7: data <= 32'hF577120C;	14'h18A8: data <= 32'hF57D2299;	14'h18A9: data <= 32'hF5833327;	14'h18AA: data <= 32'hF58943B5;	14'h18AB: data <= 32'hF58F5443;	14'h18AC: data <= 32'hF59564D1;	14'h18AD: data <= 32'hF59B755E;	14'h18AE: data <= 32'hF5A185EC;	14'h18AF: data <= 32'hF5A7967A;	14'h18B0: data <= 32'hF5ADA708;	14'h18B1: data <= 32'hF5B3B795;	14'h18B2: data <= 32'hF5B9C823;	14'h18B3: data <= 32'hF5BFD8B1;	14'h18B4: data <= 32'hF5C5E93F;	14'h18B5: data <= 32'hF5CBF9CD;	14'h18B6: data <= 32'hF5D1F717;	14'h18B7: data <= 32'hF5D7EC14;	14'h18B8: data <= 32'hF5DDE111;	14'h18B9: data <= 32'hF5E3D60E;	14'h18BA: data <= 32'hF5E9CB0B;	14'h18BB: data <= 32'hF5EFC008;	14'h18BC: data <= 32'hF5F5B505;	14'h18BD: data <= 32'hF5FBAA02;	14'h18BE: data <= 32'hF6019EFF;	14'h18BF: data <= 32'hF60793FC;	14'h18C0: data <= 32'hF60D88F8;	14'h18C1: data <= 32'hF6137DF5;	14'h18C2: data <= 32'hF61972F2;	14'h18C3: data <= 32'hF61F67EF;	14'h18C4: data <= 32'hF6255CEC;	14'h18C5: data <= 32'hF62B51E9;	14'h18C6: data <= 32'hF63146E6;	14'h18C7: data <= 32'hF6373BE3;	14'h18C8: data <= 32'hF63D30E0;	14'h18C9: data <= 32'hF64325DD;	14'h18CA: data <= 32'hF6491ADA;	14'h18CB: data <= 32'hF64F0FD7;	14'h18CC: data <= 32'hF65504D4;	14'h18CD: data <= 32'hF65AF9D1;	14'h18CE: data <= 32'hF660EECE;	14'h18CF: data <= 32'hF666E3CB;	14'h18D0: data <= 32'hF66CD8C8;	14'h18D1: data <= 32'hF672CDC5;	14'h18D2: data <= 32'hF678C2C2;	14'h18D3: data <= 32'hF67EB7BE;	14'h18D4: data <= 32'hF684ACBB;	14'h18D5: data <= 32'hF68AA1B8;	14'h18D6: data <= 32'hF69096B5;	14'h18D7: data <= 32'hF6968BB2;	14'h18D8: data <= 32'hF69C80AF;	14'h18D9: data <= 32'hF6A275AC;	14'h18DA: data <= 32'hF6A4EF1A;	14'h18DB: data <= 32'hF6A49B68;	14'h18DC: data <= 32'hF6A447B6;	14'h18DD: data <= 32'hF6A3F404;	14'h18DE: data <= 32'hF6A3A052;	14'h18DF: data <= 32'hF6A34CA0;	14'h18E0: data <= 32'hF6A2F8ED;	14'h18E1: data <= 32'hF6A2A53B;	14'h18E2: data <= 32'hF6A25189;	14'h18E3: data <= 32'hF6A1FDD7;	14'h18E4: data <= 32'hF6A1AA25;	14'h18E5: data <= 32'hF6A15673;	14'h18E6: data <= 32'hF6A102C1;	14'h18E7: data <= 32'hF6A0AF0F;	14'h18E8: data <= 32'hF6A05B5D;	14'h18E9: data <= 32'hF6A007AB;	14'h18EA: data <= 32'hF69FB3F9;	14'h18EB: data <= 32'hF69F6047;	14'h18EC: data <= 32'hF69F0C95;	14'h18ED: data <= 32'hF69EB8E3;	14'h18EE: data <= 32'hF69E6531;	14'h18EF: data <= 32'hF69E117E;	14'h18F0: data <= 32'hF69DBDCC;	14'h18F1: data <= 32'hF69D6A1A;	14'h18F2: data <= 32'hF69D1668;	14'h18F3: data <= 32'hF69CC2B6;	14'h18F4: data <= 32'hF69C6F04;	14'h18F5: data <= 32'hF69C1B52;	14'h18F6: data <= 32'hF69BC7A0;	14'h18F7: data <= 32'hF69B73EE;	14'h18F8: data <= 32'hF69B203C;	14'h18F9: data <= 32'hF69ACC8A;	14'h18FA: data <= 32'hF69A78D8;	14'h18FB: data <= 32'hF69A2526;	14'h18FC: data <= 32'hF699D174;	14'h18FD: data <= 32'hF6997DC2;	14'h18FE: data <= 32'hF697464D;	14'h18FF: data <= 32'hF69255A9;	14'h1900: data <= 32'hF68D6506;	14'h1901: data <= 32'hF6887462;	14'h1902: data <= 32'hF68383BF;	14'h1903: data <= 32'hF67E931B;	14'h1904: data <= 32'hF679A277;	14'h1905: data <= 32'hF674B1D4;	14'h1906: data <= 32'hF66FC130;	14'h1907: data <= 32'hF66AD08C;	14'h1908: data <= 32'hF665DFE9;	14'h1909: data <= 32'hF660EF45;	14'h190A: data <= 32'hF65BFEA2;	14'h190B: data <= 32'hF6570DFE;	14'h190C: data <= 32'hF6521D5A;	14'h190D: data <= 32'hF64D2CB7;	14'h190E: data <= 32'hF6483C13;	14'h190F: data <= 32'hF6434B70;	14'h1910: data <= 32'hF63E5ACC;	14'h1911: data <= 32'hF6396A28;	14'h1912: data <= 32'hF6347985;	14'h1913: data <= 32'hF62F88E1;	14'h1914: data <= 32'hF62A983D;	14'h1915: data <= 32'hF625A79A;	14'h1916: data <= 32'hF620B6F6;	14'h1917: data <= 32'hF61BC653;	14'h1918: data <= 32'hF616D5AF;	14'h1919: data <= 32'hF611E50B;	14'h191A: data <= 32'hF60CF468;	14'h191B: data <= 32'hF60803C4;	14'h191C: data <= 32'hF6031321;	14'h191D: data <= 32'hF5FE227D;	14'h191E: data <= 32'hF5F931D9;	14'h191F: data <= 32'hF5F44136;	14'h1920: data <= 32'hF5EF5092;	14'h1921: data <= 32'hF5EA5FEE;	14'h1922: data <= 32'hF5E53C04;	14'h1923: data <= 32'hF5DF89EA;	14'h1924: data <= 32'hF5D9D7D1;	14'h1925: data <= 32'hF5D425B8;	14'h1926: data <= 32'hF5CE739F;	14'h1927: data <= 32'hF5C8C186;	14'h1928: data <= 32'hF5C30F6D;	14'h1929: data <= 32'hF5BD5D54;	14'h192A: data <= 32'hF5B7AB3B;	14'h192B: data <= 32'hF5B1F921;	14'h192C: data <= 32'hF5AC4708;	14'h192D: data <= 32'hF5A694EF;	14'h192E: data <= 32'hF5A0E2D6;	14'h192F: data <= 32'hF59B30BD;	14'h1930: data <= 32'hF5957EA4;	14'h1931: data <= 32'hF58FCC8B;	14'h1932: data <= 32'hF58A1A71;	14'h1933: data <= 32'hF5846858;	14'h1934: data <= 32'hF57EB63F;	14'h1935: data <= 32'hF5790426;	14'h1936: data <= 32'hF573520D;	14'h1937: data <= 32'hF56D9FF4;	14'h1938: data <= 32'hF567EDDB;	14'h1939: data <= 32'hF5623BC2;	14'h193A: data <= 32'hF55C89A8;	14'h193B: data <= 32'hF556D78F;	14'h193C: data <= 32'hF5512576;	14'h193D: data <= 32'hF54B735D;	14'h193E: data <= 32'hF545C144;	14'h193F: data <= 32'hF5400F2B;	14'h1940: data <= 32'hF53A5D12;	14'h1941: data <= 32'hF534AAF8;	14'h1942: data <= 32'hF52EF8DF;	14'h1943: data <= 32'hF52946C6;	14'h1944: data <= 32'hF52394AD;	14'h1945: data <= 32'hF51DE294;	14'h1946: data <= 32'hF517E49C;	14'h1947: data <= 32'hF50FBCC5;	14'h1948: data <= 32'hF50794EE;	14'h1949: data <= 32'hF4FF6D17;	14'h194A: data <= 32'hF4F74541;	14'h194B: data <= 32'hF4EF1D6A;	14'h194C: data <= 32'hF4E6F593;	14'h194D: data <= 32'hF4DECDBC;	14'h194E: data <= 32'hF4D6A5E6;	14'h194F: data <= 32'hF4CE7E0F;	14'h1950: data <= 32'hF4C65638;	14'h1951: data <= 32'hF4BE2E62;	14'h1952: data <= 32'hF4B6068B;	14'h1953: data <= 32'hF4ADDEB4;	14'h1954: data <= 32'hF4A5B6DD;	14'h1955: data <= 32'hF49D8F07;	14'h1956: data <= 32'hF4956730;	14'h1957: data <= 32'hF48D3F59;	14'h1958: data <= 32'hF4851783;	14'h1959: data <= 32'hF47CEFAC;	14'h195A: data <= 32'hF474C7D5;	14'h195B: data <= 32'hF46C9FFE;	14'h195C: data <= 32'hF4647828;	14'h195D: data <= 32'hF45C5051;	14'h195E: data <= 32'hF454287A;	14'h195F: data <= 32'hF44C00A4;	14'h1960: data <= 32'hF443D8CD;	14'h1961: data <= 32'hF43BB0F6;	14'h1962: data <= 32'hF433891F;	14'h1963: data <= 32'hF42B6149;	14'h1964: data <= 32'hF4233972;	14'h1965: data <= 32'hF41B119B;	14'h1966: data <= 32'hF412E9C5;	14'h1967: data <= 32'hF40AC1EE;	14'h1968: data <= 32'hF4029A17;	14'h1969: data <= 32'hF3FA7240;	14'h196A: data <= 32'hF3F24A6A;	14'h196B: data <= 32'hF3F0D650;	14'h196C: data <= 32'hF3EF8C94;	14'h196D: data <= 32'hF3EE42D8;	14'h196E: data <= 32'hF3ECF91C;	14'h196F: data <= 32'hF3EBAF60;	14'h1970: data <= 32'hF3EA65A4;	14'h1971: data <= 32'hF3E91BE8;	14'h1972: data <= 32'hF3E7D22C;	14'h1973: data <= 32'hF3E68870;	14'h1974: data <= 32'hF3E53EB4;	14'h1975: data <= 32'hF3E3F4F8;	14'h1976: data <= 32'hF3E2AB3C;	14'h1977: data <= 32'hF3E16180;	14'h1978: data <= 32'hF3E017C4;	14'h1979: data <= 32'hF3DECE08;	14'h197A: data <= 32'hF3DD844C;	14'h197B: data <= 32'hF3DC3A90;	14'h197C: data <= 32'hF3DAF0D4;	14'h197D: data <= 32'hF3D9A718;	14'h197E: data <= 32'hF3D85D5B;	14'h197F: data <= 32'hF3D7139F;	14'h1980: data <= 32'hF3D5C9E3;	14'h1981: data <= 32'hF3D48027;	14'h1982: data <= 32'hF3D3366B;	14'h1983: data <= 32'hF3D1ECAF;	14'h1984: data <= 32'hF3D0A2F3;	14'h1985: data <= 32'hF3CF5937;	14'h1986: data <= 32'hF3CE0F7B;	14'h1987: data <= 32'hF3CCC5BF;	14'h1988: data <= 32'hF3CB7C03;	14'h1989: data <= 32'hF3CA3247;	14'h198A: data <= 32'hF3C8E88B;	14'h198B: data <= 32'hF3C79ECF;	14'h198C: data <= 32'hF3C65513;	14'h198D: data <= 32'hF3C50B57;	14'h198E: data <= 32'hF3C3C19B;	14'h198F: data <= 32'hF3C2D18D;	14'h1990: data <= 32'hF3C1F3B2;	14'h1991: data <= 32'hF3C115D6;	14'h1992: data <= 32'hF3C037FB;	14'h1993: data <= 32'hF3BF5A20;	14'h1994: data <= 32'hF3BE7C44;	14'h1995: data <= 32'hF3BD9E69;	14'h1996: data <= 32'hF3BCC08E;	14'h1997: data <= 32'hF3BBE2B2;	14'h1998: data <= 32'hF3BB04D7;	14'h1999: data <= 32'hF3BA26FC;	14'h199A: data <= 32'hF3B94920;	14'h199B: data <= 32'hF3B86B45;	14'h199C: data <= 32'hF3B78D6A;	14'h199D: data <= 32'hF3B6AF8E;	14'h199E: data <= 32'hF3B5D1B3;	14'h199F: data <= 32'hF3B4F3D7;	14'h19A0: data <= 32'hF3B415FC;	14'h19A1: data <= 32'hF3B33821;	14'h19A2: data <= 32'hF3B25A45;	14'h19A3: data <= 32'hF3B17C6A;	14'h19A4: data <= 32'hF3B09E8F;	14'h19A5: data <= 32'hF3AFC0B3;	14'h19A6: data <= 32'hF3AEE2D8;	14'h19A7: data <= 32'hF3AE04FD;	14'h19A8: data <= 32'hF3AD2721;	14'h19A9: data <= 32'hF3AC4946;	14'h19AA: data <= 32'hF3AB6B6B;	14'h19AB: data <= 32'hF3AA8D8F;	14'h19AC: data <= 32'hF3A9AFB4;	14'h19AD: data <= 32'hF3A8D1D9;	14'h19AE: data <= 32'hF3A7F3FD;	14'h19AF: data <= 32'hF3A71622;	14'h19B0: data <= 32'hF3A63847;	14'h19B1: data <= 32'hF3A55A6B;	14'h19B2: data <= 32'hF3A47C90;	14'h19B3: data <= 32'hF3A495C2;	14'h19B4: data <= 32'hF3A51FA4;	14'h19B5: data <= 32'hF3A5A986;	14'h19B6: data <= 32'hF3A63368;	14'h19B7: data <= 32'hF3A6BD4B;	14'h19B8: data <= 32'hF3A7472D;	14'h19B9: data <= 32'hF3A7D10F;	14'h19BA: data <= 32'hF3A85AF2;	14'h19BB: data <= 32'hF3A8E4D4;	14'h19BC: data <= 32'hF3A96EB6;	14'h19BD: data <= 32'hF3A9F899;	14'h19BE: data <= 32'hF3AA827B;	14'h19BF: data <= 32'hF3AB0C5D;	14'h19C0: data <= 32'hF3AB9640;	14'h19C1: data <= 32'hF3AC2022;	14'h19C2: data <= 32'hF3ACAA04;	14'h19C3: data <= 32'hF3AD33E7;	14'h19C4: data <= 32'hF3ADBDC9;	14'h19C5: data <= 32'hF3AE47AB;	14'h19C6: data <= 32'hF3AED18E;	14'h19C7: data <= 32'hF3AF5B70;	14'h19C8: data <= 32'hF3AFE552;	14'h19C9: data <= 32'hF3B06F35;	14'h19CA: data <= 32'hF3B0F917;	14'h19CB: data <= 32'hF3B182F9;	14'h19CC: data <= 32'hF3B20CDC;	14'h19CD: data <= 32'hF3B296BE;	14'h19CE: data <= 32'hF3B320A0;	14'h19CF: data <= 32'hF3B3AA83;	14'h19D0: data <= 32'hF3B43465;	14'h19D1: data <= 32'hF3B4BE47;	14'h19D2: data <= 32'hF3B5482A;	14'h19D3: data <= 32'hF3B5D20C;	14'h19D4: data <= 32'hF3B65BEE;	14'h19D5: data <= 32'hF3B6E5D0;	14'h19D6: data <= 32'hF3B76FB3;	14'h19D7: data <= 32'hF3B8EE54;	14'h19D8: data <= 32'hF3BB3BA3;	14'h19D9: data <= 32'hF3BD88F2;	14'h19DA: data <= 32'hF3BFD640;	14'h19DB: data <= 32'hF3C2238F;	14'h19DC: data <= 32'hF3C470DD;	14'h19DD: data <= 32'hF3C6BE2C;	14'h19DE: data <= 32'hF3C90B7B;	14'h19DF: data <= 32'hF3CB58C9;	14'h19E0: data <= 32'hF3CDA618;	14'h19E1: data <= 32'hF3CFF366;	14'h19E2: data <= 32'hF3D240B5;	14'h19E3: data <= 32'hF3D48E04;	14'h19E4: data <= 32'hF3D6DB52;	14'h19E5: data <= 32'hF3D928A1;	14'h19E6: data <= 32'hF3DB75EF;	14'h19E7: data <= 32'hF3DDC33E;	14'h19E8: data <= 32'hF3E0108D;	14'h19E9: data <= 32'hF3E25DDB;	14'h19EA: data <= 32'hF3E4AB2A;	14'h19EB: data <= 32'hF3E6F878;	14'h19EC: data <= 32'hF3E945C7;	14'h19ED: data <= 32'hF3EB9316;	14'h19EE: data <= 32'hF3EDE064;	14'h19EF: data <= 32'hF3F02DB3;	14'h19F0: data <= 32'hF3F27B01;	14'h19F1: data <= 32'hF3F4C850;	14'h19F2: data <= 32'hF3F7159F;	14'h19F3: data <= 32'hF3F962ED;	14'h19F4: data <= 32'hF3FBB03C;	14'h19F5: data <= 32'hF3FDFD8A;	14'h19F6: data <= 32'hF4004AD9;	14'h19F7: data <= 32'hF4029828;	14'h19F8: data <= 32'hF404E576;	14'h19F9: data <= 32'hF40732C5;	14'h19FA: data <= 32'hF4098013;	14'h19FB: data <= 32'hF40AC5B5;	14'h19FC: data <= 32'hF40A7BD4;	14'h19FD: data <= 32'hF40A31F3;	14'h19FE: data <= 32'hF409E812;	14'h19FF: data <= 32'hF4099E32;	14'h1A00: data <= 32'hF4095451;	14'h1A01: data <= 32'hF4090A70;	14'h1A02: data <= 32'hF408C08F;	14'h1A03: data <= 32'hF40876AE;	14'h1A04: data <= 32'hF4082CCD;	14'h1A05: data <= 32'hF407E2EC;	14'h1A06: data <= 32'hF407990C;	14'h1A07: data <= 32'hF4074F2B;	14'h1A08: data <= 32'hF407054A;	14'h1A09: data <= 32'hF406BB69;	14'h1A0A: data <= 32'hF4067188;	14'h1A0B: data <= 32'hF40627A7;	14'h1A0C: data <= 32'hF405DDC6;	14'h1A0D: data <= 32'hF40593E6;	14'h1A0E: data <= 32'hF4054A05;	14'h1A0F: data <= 32'hF4050024;	14'h1A10: data <= 32'hF404B643;	14'h1A11: data <= 32'hF4046C62;	14'h1A12: data <= 32'hF4042281;	14'h1A13: data <= 32'hF403D8A1;	14'h1A14: data <= 32'hF4038EC0;	14'h1A15: data <= 32'hF40344DF;	14'h1A16: data <= 32'hF402FAFE;	14'h1A17: data <= 32'hF402B11D;	14'h1A18: data <= 32'hF402673C;	14'h1A19: data <= 32'hF4021D5B;	14'h1A1A: data <= 32'hF401D37B;	14'h1A1B: data <= 32'hF401899A;	14'h1A1C: data <= 32'hF4013FB9;	14'h1A1D: data <= 32'hF400F5D8;	14'h1A1E: data <= 32'hF400ABF7;	14'h1A1F: data <= 32'hF3FE90DD;	14'h1A20: data <= 32'hF3F7183C;	14'h1A21: data <= 32'hF3EF9F9B;	14'h1A22: data <= 32'hF3E826FB;	14'h1A23: data <= 32'hF3E0AE5A;	14'h1A24: data <= 32'hF3D935BA;	14'h1A25: data <= 32'hF3D1BD19;	14'h1A26: data <= 32'hF3CA4479;	14'h1A27: data <= 32'hF3C2CBD8;	14'h1A28: data <= 32'hF3BB5337;	14'h1A29: data <= 32'hF3B3DA97;	14'h1A2A: data <= 32'hF3AC61F6;	14'h1A2B: data <= 32'hF3A4E956;	14'h1A2C: data <= 32'hF39D70B5;	14'h1A2D: data <= 32'hF395F814;	14'h1A2E: data <= 32'hF38E7F74;	14'h1A2F: data <= 32'hF38706D3;	14'h1A30: data <= 32'hF37F8E33;	14'h1A31: data <= 32'hF3781592;	14'h1A32: data <= 32'hF3709CF2;	14'h1A33: data <= 32'hF3692451;	14'h1A34: data <= 32'hF361ABB0;	14'h1A35: data <= 32'hF35A3310;	14'h1A36: data <= 32'hF352BA6F;	14'h1A37: data <= 32'hF34B41CF;	14'h1A38: data <= 32'hF343C92E;	14'h1A39: data <= 32'hF33C508E;	14'h1A3A: data <= 32'hF334D7ED;	14'h1A3B: data <= 32'hF32D5F4C;	14'h1A3C: data <= 32'hF325E6AC;	14'h1A3D: data <= 32'hF31E6E0B;	14'h1A3E: data <= 32'hF316F56B;	14'h1A3F: data <= 32'hF30F7CCA;	14'h1A40: data <= 32'hF308042A;	14'h1A41: data <= 32'hF3008B89;	14'h1A42: data <= 32'hF2F912E8;	14'h1A43: data <= 32'hF2F0CC1F;	14'h1A44: data <= 32'hF2E1E63C;	14'h1A45: data <= 32'hF2D3005A;	14'h1A46: data <= 32'hF2C41A77;	14'h1A47: data <= 32'hF2B53495;	14'h1A48: data <= 32'hF2A64EB3;	14'h1A49: data <= 32'hF29768D0;	14'h1A4A: data <= 32'hF28882EE;	14'h1A4B: data <= 32'hF2799D0B;	14'h1A4C: data <= 32'hF26AB729;	14'h1A4D: data <= 32'hF25BD146;	14'h1A4E: data <= 32'hF24CEB64;	14'h1A4F: data <= 32'hF23E0582;	14'h1A50: data <= 32'hF22F1F9F;	14'h1A51: data <= 32'hF22039BD;	14'h1A52: data <= 32'hF21153DA;	14'h1A53: data <= 32'hF2026DF8;	14'h1A54: data <= 32'hF1F38816;	14'h1A55: data <= 32'hF1E4A233;	14'h1A56: data <= 32'hF1D5BC51;	14'h1A57: data <= 32'hF1C6D66E;	14'h1A58: data <= 32'hF1B7F08C;	14'h1A59: data <= 32'hF1A90AA9;	14'h1A5A: data <= 32'hF19A24C7;	14'h1A5B: data <= 32'hF18B3EE5;	14'h1A5C: data <= 32'hF17C5902;	14'h1A5D: data <= 32'hF16D7320;	14'h1A5E: data <= 32'hF15E8D3D;	14'h1A5F: data <= 32'hF14FA75B;	14'h1A60: data <= 32'hF140C178;	14'h1A61: data <= 32'hF131DB96;	14'h1A62: data <= 32'hF122F5B4;	14'h1A63: data <= 32'hF1140FD1;	14'h1A64: data <= 32'hF10529EF;	14'h1A65: data <= 32'hF0F6440C;	14'h1A66: data <= 32'hF0E75E2A;	14'h1A67: data <= 32'hF0D87847;	14'h1A68: data <= 32'hF0C20457;	14'h1A69: data <= 32'hF0AB47DF;	14'h1A6A: data <= 32'hF0948B67;	14'h1A6B: data <= 32'hF07DCEEF;	14'h1A6C: data <= 32'hF0671277;	14'h1A6D: data <= 32'hF05055FF;	14'h1A6E: data <= 32'hF0399988;	14'h1A6F: data <= 32'hF022DD10;	14'h1A70: data <= 32'hF00C2098;	14'h1A71: data <= 32'hEFF56420;	14'h1A72: data <= 32'hEFDEA7A8;	14'h1A73: data <= 32'hEFC7EB31;	14'h1A74: data <= 32'hEFB12EB9;	14'h1A75: data <= 32'hEF9A7241;	14'h1A76: data <= 32'hEF83B5C9;	14'h1A77: data <= 32'hEF6CF951;	14'h1A78: data <= 32'hEF563CD9;	14'h1A79: data <= 32'hEF3F8062;	14'h1A7A: data <= 32'hEF28C3EA;	14'h1A7B: data <= 32'hEF120772;	14'h1A7C: data <= 32'hEEFB4AFA;	14'h1A7D: data <= 32'hEEE48E82;	14'h1A7E: data <= 32'hEECDD20A;	14'h1A7F: data <= 32'hEEB71593;	14'h1A80: data <= 32'hEEA0591B;	14'h1A81: data <= 32'hEE899CA3;	14'h1A82: data <= 32'hEE72E02B;	14'h1A83: data <= 32'hEE5C23B3;	14'h1A84: data <= 32'hEE45673C;	14'h1A85: data <= 32'hEE2EAAC4;	14'h1A86: data <= 32'hEE17EE4C;	14'h1A87: data <= 32'hEE0131D4;	14'h1A88: data <= 32'hEDEA755C;	14'h1A89: data <= 32'hEDD3B8E4;	14'h1A8A: data <= 32'hEDBCFC6D;	14'h1A8B: data <= 32'hEDA63FF5;	14'h1A8C: data <= 32'hED8E47C4;	14'h1A8D: data <= 32'hED7609EF;	14'h1A8E: data <= 32'hED5DCC1A;	14'h1A8F: data <= 32'hED458E44;	14'h1A90: data <= 32'hED2D506F;	14'h1A91: data <= 32'hED15129A;	14'h1A92: data <= 32'hECFCD4C4;	14'h1A93: data <= 32'hECE496EF;	14'h1A94: data <= 32'hECCC591A;	14'h1A95: data <= 32'hECB41B44;	14'h1A96: data <= 32'hEC9BDD6F;	14'h1A97: data <= 32'hEC839F9A;	14'h1A98: data <= 32'hEC6B61C4;	14'h1A99: data <= 32'hEC5323EF;	14'h1A9A: data <= 32'hEC3AE61A;	14'h1A9B: data <= 32'hEC22A844;	14'h1A9C: data <= 32'hEC0A6A6F;	14'h1A9D: data <= 32'hEBF22C9A;	14'h1A9E: data <= 32'hEBD9EEC4;	14'h1A9F: data <= 32'hEBC1B0EF;	14'h1AA0: data <= 32'hEBA9731A;	14'h1AA1: data <= 32'hEB913544;	14'h1AA2: data <= 32'hEB78F76F;	14'h1AA3: data <= 32'hEB60B999;	14'h1AA4: data <= 32'hEB487BC4;	14'h1AA5: data <= 32'hEB303DEF;	14'h1AA6: data <= 32'hEB180019;	14'h1AA7: data <= 32'hEAFFC244;	14'h1AA8: data <= 32'hEAE7846F;	14'h1AA9: data <= 32'hEACF4699;	14'h1AAA: data <= 32'hEAB708C4;	14'h1AAB: data <= 32'hEA9ECAEF;	14'h1AAC: data <= 32'hEA868D19;	14'h1AAD: data <= 32'hEA6E4F44;	14'h1AAE: data <= 32'hEA56116F;	14'h1AAF: data <= 32'hEA3DD399;	14'h1AB0: data <= 32'hEA29530C;	14'h1AB1: data <= 32'hEA16A00B;	14'h1AB2: data <= 32'hEA03ED0A;	14'h1AB3: data <= 32'hE9F13A0A;	14'h1AB4: data <= 32'hE9DE8709;	14'h1AB5: data <= 32'hE9CBD408;	14'h1AB6: data <= 32'hE9B92107;	14'h1AB7: data <= 32'hE9A66E06;	14'h1AB8: data <= 32'hE993BB05;	14'h1AB9: data <= 32'hE9810804;	14'h1ABA: data <= 32'hE96E5503;	14'h1ABB: data <= 32'hE95BA202;	14'h1ABC: data <= 32'hE948EF01;	14'h1ABD: data <= 32'hE9363C00;	14'h1ABE: data <= 32'hE92388FF;	14'h1ABF: data <= 32'hE910D5FE;	14'h1AC0: data <= 32'hE8FE22FD;	14'h1AC1: data <= 32'hE8EB6FFC;	14'h1AC2: data <= 32'hE8D8BCFB;	14'h1AC3: data <= 32'hE8C609FA;	14'h1AC4: data <= 32'hE8B356F9;	14'h1AC5: data <= 32'hE8A0A3F8;	14'h1AC6: data <= 32'hE88DF0F7;	14'h1AC7: data <= 32'hE87B3DF7;	14'h1AC8: data <= 32'hE8688AF6;	14'h1AC9: data <= 32'hE855D7F5;	14'h1ACA: data <= 32'hE84324F4;	14'h1ACB: data <= 32'hE83071F3;	14'h1ACC: data <= 32'hE81DBEF2;	14'h1ACD: data <= 32'hE80B0BF1;	14'h1ACE: data <= 32'hE7F858F0;	14'h1ACF: data <= 32'hE7E5A5EF;	14'h1AD0: data <= 32'hE7D2F2EE;	14'h1AD1: data <= 32'hE7C03FED;	14'h1AD2: data <= 32'hE7AD8CEC;	14'h1AD3: data <= 32'hE79AD9EB;	14'h1AD4: data <= 32'hE7894A9E;	14'h1AD5: data <= 32'hE778BDE0;	14'h1AD6: data <= 32'hE7683122;	14'h1AD7: data <= 32'hE757A464;	14'h1AD8: data <= 32'hE74717A5;	14'h1AD9: data <= 32'hE7368AE7;	14'h1ADA: data <= 32'hE725FE29;	14'h1ADB: data <= 32'hE715716A;	14'h1ADC: data <= 32'hE704E4AC;	14'h1ADD: data <= 32'hE6F457EE;	14'h1ADE: data <= 32'hE6E3CB2F;	14'h1ADF: data <= 32'hE6D33E71;	14'h1AE0: data <= 32'hE6C2B1B3;	14'h1AE1: data <= 32'hE6B224F4;	14'h1AE2: data <= 32'hE6A19836;	14'h1AE3: data <= 32'hE6910B78;	14'h1AE4: data <= 32'hE6807EB9;	14'h1AE5: data <= 32'hE66FF1FB;	14'h1AE6: data <= 32'hE65F653D;	14'h1AE7: data <= 32'hE64ED87E;	14'h1AE8: data <= 32'hE63E4BC0;	14'h1AE9: data <= 32'hE62DBF02;	14'h1AEA: data <= 32'hE61D3243;	14'h1AEB: data <= 32'hE60CA585;	14'h1AEC: data <= 32'hE5FC18C7;	14'h1AED: data <= 32'hE5EB8C09;	14'h1AEE: data <= 32'hE5DAFF4A;	14'h1AEF: data <= 32'hE5CA728C;	14'h1AF0: data <= 32'hE5B9E5CE;	14'h1AF1: data <= 32'hE5A9590F;	14'h1AF2: data <= 32'hE598CC51;	14'h1AF3: data <= 32'hE5883F93;	14'h1AF4: data <= 32'hE577B2D4;	14'h1AF5: data <= 32'hE5672616;	14'h1AF6: data <= 32'hE5569958;	14'h1AF7: data <= 32'hE5460C99;	14'h1AF8: data <= 32'hE53273F8;	14'h1AF9: data <= 32'hE51A0064;	14'h1AFA: data <= 32'hE5018CD0;	14'h1AFB: data <= 32'hE4E9193C;	14'h1AFC: data <= 32'hE4D0A5A8;	14'h1AFD: data <= 32'hE4B83214;	14'h1AFE: data <= 32'hE49FBE80;	14'h1AFF: data <= 32'hE4874AEC;	14'h1B00: data <= 32'hE46ED758;	14'h1B01: data <= 32'hE45663C4;	14'h1B02: data <= 32'hE43DF030;	14'h1B03: data <= 32'hE4257C9C;	14'h1B04: data <= 32'hE40D0908;	14'h1B05: data <= 32'hE3F49574;	14'h1B06: data <= 32'hE3DC21E0;	14'h1B07: data <= 32'hE3C3AE4C;	14'h1B08: data <= 32'hE3AB3AB8;	14'h1B09: data <= 32'hE392C724;	14'h1B0A: data <= 32'hE37A5390;	14'h1B0B: data <= 32'hE361DFFC;	14'h1B0C: data <= 32'hE3496C68;	14'h1B0D: data <= 32'hE330F8D4;	14'h1B0E: data <= 32'hE3188540;	14'h1B0F: data <= 32'hE30011AC;	14'h1B10: data <= 32'hE2E79E18;	14'h1B11: data <= 32'hE2CF2A84;	14'h1B12: data <= 32'hE2B6B6F0;	14'h1B13: data <= 32'hE29E435C;	14'h1B14: data <= 32'hE285CFC8;	14'h1B15: data <= 32'hE26D5C34;	14'h1B16: data <= 32'hE254E8A0;	14'h1B17: data <= 32'hE23C750C;	14'h1B18: data <= 32'hE2240178;	14'h1B19: data <= 32'hE20B8DE4;	14'h1B1A: data <= 32'hE1F31A4F;	14'h1B1B: data <= 32'hE1DAA6BB;	14'h1B1C: data <= 32'hE1C0D319;	14'h1B1D: data <= 32'hE1A2AA7B;	14'h1B1E: data <= 32'hE18481DD;	14'h1B1F: data <= 32'hE1665940;	14'h1B20: data <= 32'hE14830A2;	14'h1B21: data <= 32'hE12A0804;	14'h1B22: data <= 32'hE10BDF67;	14'h1B23: data <= 32'hE0EDB6C9;	14'h1B24: data <= 32'hE0CF8E2B;	14'h1B25: data <= 32'hE0B1658E;	14'h1B26: data <= 32'hE0933CF0;	14'h1B27: data <= 32'hE0751452;	14'h1B28: data <= 32'hE056EBB5;	14'h1B29: data <= 32'hE038C317;	14'h1B2A: data <= 32'hE01A9A79;	14'h1B2B: data <= 32'hDFFC71DC;	14'h1B2C: data <= 32'hDFDE493E;	14'h1B2D: data <= 32'hDFC020A0;	14'h1B2E: data <= 32'hDFA1F803;	14'h1B2F: data <= 32'hDF83CF65;	14'h1B30: data <= 32'hDF65A6C7;	14'h1B31: data <= 32'hDF477E2A;	14'h1B32: data <= 32'hDF29558C;	14'h1B33: data <= 32'hDF0B2CEE;	14'h1B34: data <= 32'hDEED0451;	14'h1B35: data <= 32'hDECEDBB3;	14'h1B36: data <= 32'hDEB0B315;	14'h1B37: data <= 32'hDE928A78;	14'h1B38: data <= 32'hDE7461DA;	14'h1B39: data <= 32'hDE56393C;	14'h1B3A: data <= 32'hDE38109F;	14'h1B3B: data <= 32'hDE19E801;	14'h1B3C: data <= 32'hDDFBBF63;	14'h1B3D: data <= 32'hDDDD96C6;	14'h1B3E: data <= 32'hDDBF6E28;	14'h1B3F: data <= 32'hDDA1458A;	14'h1B40: data <= 32'hDD8256E5;	14'h1B41: data <= 32'hDD5C27B8;	14'h1B42: data <= 32'hDD35F88B;	14'h1B43: data <= 32'hDD0FC95E;	14'h1B44: data <= 32'hDCE99A31;	14'h1B45: data <= 32'hDCC36B03;	14'h1B46: data <= 32'hDC9D3BD6;	14'h1B47: data <= 32'hDC770CA9;	14'h1B48: data <= 32'hDC50DD7C;	14'h1B49: data <= 32'hDC2AAE4F;	14'h1B4A: data <= 32'hDC047F22;	14'h1B4B: data <= 32'hDBDE4FF5;	14'h1B4C: data <= 32'hDBB820C8;	14'h1B4D: data <= 32'hDB91F19B;	14'h1B4E: data <= 32'hDB6BC26E;	14'h1B4F: data <= 32'hDB459340;	14'h1B50: data <= 32'hDB1F6413;	14'h1B51: data <= 32'hDAF934E6;	14'h1B52: data <= 32'hDAD305B9;	14'h1B53: data <= 32'hDAACD68C;	14'h1B54: data <= 32'hDA86A75F;	14'h1B55: data <= 32'hDA607832;	14'h1B56: data <= 32'hDA3A4905;	14'h1B57: data <= 32'hDA1419D8;	14'h1B58: data <= 32'hD9EDEAAA;	14'h1B59: data <= 32'hD9C7BB7D;	14'h1B5A: data <= 32'hD9A18C50;	14'h1B5B: data <= 32'hD97B5D23;	14'h1B5C: data <= 32'hD9552DF6;	14'h1B5D: data <= 32'hD92EFEC9;	14'h1B5E: data <= 32'hD908CF9C;	14'h1B5F: data <= 32'hD8E2A06F;	14'h1B60: data <= 32'hD8BC7142;	14'h1B61: data <= 32'hD8964215;	14'h1B62: data <= 32'hD87012E7;	14'h1B63: data <= 32'hD849E3BA;	14'h1B64: data <= 32'hD823B48D;	14'h1B65: data <= 32'hD7ED9DB2;	14'h1B66: data <= 32'hD7B6B8AD;	14'h1B67: data <= 32'hD77FD3A8;	14'h1B68: data <= 32'hD748EEA4;	14'h1B69: data <= 32'hD712099F;	14'h1B6A: data <= 32'hD6DB249A;	14'h1B6B: data <= 32'hD6A43F95;	14'h1B6C: data <= 32'hD66D5A91;	14'h1B6D: data <= 32'hD636758C;	14'h1B6E: data <= 32'hD5FF9087;	14'h1B6F: data <= 32'hD5C8AB82;	14'h1B70: data <= 32'hD591C67E;	14'h1B71: data <= 32'hD55AE179;	14'h1B72: data <= 32'hD523FC74;	14'h1B73: data <= 32'hD4ED176F;	14'h1B74: data <= 32'hD4B6326A;	14'h1B75: data <= 32'hD47F4D66;	14'h1B76: data <= 32'hD4486861;	14'h1B77: data <= 32'hD411835C;	14'h1B78: data <= 32'hD3DA9E57;	14'h1B79: data <= 32'hD3A3B953;	14'h1B7A: data <= 32'hD36CD44E;	14'h1B7B: data <= 32'hD335EF49;	14'h1B7C: data <= 32'hD2FF0A44;	14'h1B7D: data <= 32'hD2C82540;	14'h1B7E: data <= 32'hD291403B;	14'h1B7F: data <= 32'hD25A5B36;	14'h1B80: data <= 32'hD2237631;	14'h1B81: data <= 32'hD1EC912D;	14'h1B82: data <= 32'hD1B5AC28;	14'h1B83: data <= 32'hD17EC723;	14'h1B84: data <= 32'hD147E21E;	14'h1B85: data <= 32'hD110FD1A;	14'h1B86: data <= 32'hD0DA1815;	14'h1B87: data <= 32'hD0A33310;	14'h1B88: data <= 32'hD06C4E0B;	14'h1B89: data <= 32'hD0255227;	14'h1B8A: data <= 32'hCFDA7EA7;	14'h1B8B: data <= 32'hCF8FAB26;	14'h1B8C: data <= 32'hCF44D7A5;	14'h1B8D: data <= 32'hCEFA0425;	14'h1B8E: data <= 32'hCEAF30A4;	14'h1B8F: data <= 32'hCE645D23;	14'h1B90: data <= 32'hCE1989A3;	14'h1B91: data <= 32'hCDCEB622;	14'h1B92: data <= 32'hCD83E2A1;	14'h1B93: data <= 32'hCD390F21;	14'h1B94: data <= 32'hCCEE3BA0;	14'h1B95: data <= 32'hCCA3681F;	14'h1B96: data <= 32'hCC58949F;	14'h1B97: data <= 32'hCC0DC11E;	14'h1B98: data <= 32'hCBC2ED9E;	14'h1B99: data <= 32'hCB781A1D;	14'h1B9A: data <= 32'hCB2D469C;	14'h1B9B: data <= 32'hCAE2731C;	14'h1B9C: data <= 32'hCA979F9B;	14'h1B9D: data <= 32'hCA4CCC1A;	14'h1B9E: data <= 32'hCA01F89A;	14'h1B9F: data <= 32'hC9B72519;	14'h1BA0: data <= 32'hC96C5198;	14'h1BA1: data <= 32'hC9217E18;	14'h1BA2: data <= 32'hC8D6AA97;	14'h1BA3: data <= 32'hC88BD716;	14'h1BA4: data <= 32'hC8410396;	14'h1BA5: data <= 32'hC7F63015;	14'h1BA6: data <= 32'hC7AB5C94;	14'h1BA7: data <= 32'hC7608914;	14'h1BA8: data <= 32'hC715B593;	14'h1BA9: data <= 32'hC6CAE212;	14'h1BAA: data <= 32'hC6800E92;	14'h1BAB: data <= 32'hC6353B11;	14'h1BAC: data <= 32'hC5EA6790;	14'h1BAD: data <= 32'hC57A6295;	14'h1BAE: data <= 32'hC4F76E4E;	14'h1BAF: data <= 32'hC4747A07;	14'h1BB0: data <= 32'hC3F185BF;	14'h1BB1: data <= 32'hC36E9178;	14'h1BB2: data <= 32'hC2EB9D30;	14'h1BB3: data <= 32'hC268A8E9;	14'h1BB4: data <= 32'hC1E5B4A2;	14'h1BB5: data <= 32'hC162C05A;	14'h1BB6: data <= 32'hC0DFCC13;	14'h1BB7: data <= 32'hC05CD7CB;	14'h1BB8: data <= 32'hBFD9E384;	14'h1BB9: data <= 32'hBF56EF3D;	14'h1BBA: data <= 32'hBED3FAF5;	14'h1BBB: data <= 32'hBE5106AE;	14'h1BBC: data <= 32'hBDCE1267;	14'h1BBD: data <= 32'hBD4B1E1F;	14'h1BBE: data <= 32'hBCC829D8;	14'h1BBF: data <= 32'hBC453590;	14'h1BC0: data <= 32'hBBC24149;	14'h1BC1: data <= 32'hBB3F4D02;	14'h1BC2: data <= 32'hBABC58BA;	14'h1BC3: data <= 32'hBA396473;	14'h1BC4: data <= 32'hB9B6702C;	14'h1BC5: data <= 32'hB9337BE4;	14'h1BC6: data <= 32'hB8B0879D;	14'h1BC7: data <= 32'hB82D9355;	14'h1BC8: data <= 32'hB7AA9F0E;	14'h1BC9: data <= 32'hB727AAC7;	14'h1BCA: data <= 32'hB6A4B67F;	14'h1BCB: data <= 32'hB621C238;	14'h1BCC: data <= 32'hB59ECDF0;	14'h1BCD: data <= 32'hB51BD9A9;	14'h1BCE: data <= 32'hB498E562;	14'h1BCF: data <= 32'hB415F11A;	14'h1BD0: data <= 32'hB392FCD3;	14'h1BD1: data <= 32'hB29789F5;	14'h1BD2: data <= 32'hB12C0096;	14'h1BD3: data <= 32'hAFC07738;	14'h1BD4: data <= 32'hAE54EDD9;	14'h1BD5: data <= 32'hACE9647A;	14'h1BD6: data <= 32'hAB7DDB1C;	14'h1BD7: data <= 32'hAA1251BD;	14'h1BD8: data <= 32'hA8A6C85F;	14'h1BD9: data <= 32'hA73B3F00;	14'h1BDA: data <= 32'hA5CFB5A1;	14'h1BDB: data <= 32'hA4642C43;	14'h1BDC: data <= 32'hA2F8A2E4;	14'h1BDD: data <= 32'hA18D1986;	14'h1BDE: data <= 32'hA0219027;	14'h1BDF: data <= 32'h9EB606C9;	14'h1BE0: data <= 32'h9D4A7D6A;	14'h1BE1: data <= 32'h9BDEF40B;	14'h1BE2: data <= 32'h9A736AAD;	14'h1BE3: data <= 32'h9907E14E;	14'h1BE4: data <= 32'h979C57F0;	14'h1BE5: data <= 32'h9630CE91;	14'h1BE6: data <= 32'h94C54532;	14'h1BE7: data <= 32'h9359BBD4;	14'h1BE8: data <= 32'h91EE3275;	14'h1BE9: data <= 32'h9082A917;	14'h1BEA: data <= 32'h8F171FB8;	14'h1BEB: data <= 32'h8DAB965A;	14'h1BEC: data <= 32'h8C400CFB;	14'h1BED: data <= 32'h8AD4839C;	14'h1BEE: data <= 32'h8968FA3E;	14'h1BEF: data <= 32'h87FD70DF;	14'h1BF0: data <= 32'h8691E781;	14'h1BF1: data <= 32'h85265E22;	14'h1BF2: data <= 32'h83BAD4C3;	14'h1BF3: data <= 32'h824F4B65;	14'h1BF4: data <= 32'h80E3C206;	14'h1BF5: data <= 32'h809149F5;	14'h1BF6: data <= 32'h821649C2;	14'h1BF7: data <= 32'h839B498E;	14'h1BF8: data <= 32'h8520495B;	14'h1BF9: data <= 32'h86A54928;	14'h1BFA: data <= 32'h882A48F4;	14'h1BFB: data <= 32'h89AF48C1;	14'h1BFC: data <= 32'h8B34488D;	14'h1BFD: data <= 32'h8CB9485A;	14'h1BFE: data <= 32'h8E3E4826;	14'h1BFF: data <= 32'h8FC347F3;	14'h1C00: data <= 32'h914847BF;	14'h1C01: data <= 32'h92CD478C;	14'h1C02: data <= 32'h94524758;	14'h1C03: data <= 32'h95D74725;	14'h1C04: data <= 32'h975C46F1;	14'h1C05: data <= 32'h98E146BE;	14'h1C06: data <= 32'h9A66468A;	14'h1C07: data <= 32'h9BEB4657;	14'h1C08: data <= 32'h9D704623;	14'h1C09: data <= 32'h9EF545F0;	14'h1C0A: data <= 32'hA07A45BC;	14'h1C0B: data <= 32'hA1FF4589;	14'h1C0C: data <= 32'hA3844555;	14'h1C0D: data <= 32'hA5094522;	14'h1C0E: data <= 32'hA68E44EE;	14'h1C0F: data <= 32'hA81344BB;	14'h1C10: data <= 32'hA9984487;	14'h1C11: data <= 32'hAB1D4454;	14'h1C12: data <= 32'hACA24420;	14'h1C13: data <= 32'hAE2743ED;	14'h1C14: data <= 32'hAFAC43B9;	14'h1C15: data <= 32'hB1314386;	14'h1C16: data <= 32'hB2B64353;	14'h1C17: data <= 32'hB43B431F;	14'h1C18: data <= 32'hB5C042EC;	14'h1C19: data <= 32'hB6FE744C;	14'h1C1A: data <= 32'hB74E2440;	14'h1C1B: data <= 32'hB79DD434;	14'h1C1C: data <= 32'hB7ED8428;	14'h1C1D: data <= 32'hB83D341C;	14'h1C1E: data <= 32'hB88CE40F;	14'h1C1F: data <= 32'hB8DC9403;	14'h1C20: data <= 32'hB92C43F7;	14'h1C21: data <= 32'hB97BF3EB;	14'h1C22: data <= 32'hB9CBA3DF;	14'h1C23: data <= 32'hBA1B53D3;	14'h1C24: data <= 32'hBA6B03C7;	14'h1C25: data <= 32'hBABAB3BB;	14'h1C26: data <= 32'hBB0A63AF;	14'h1C27: data <= 32'hBB5A13A3;	14'h1C28: data <= 32'hBBA9C397;	14'h1C29: data <= 32'hBBF9738B;	14'h1C2A: data <= 32'hBC49237E;	14'h1C2B: data <= 32'hBC98D372;	14'h1C2C: data <= 32'hBCE88366;	14'h1C2D: data <= 32'hBD38335A;	14'h1C2E: data <= 32'hBD87E34E;	14'h1C2F: data <= 32'hBDD79342;	14'h1C30: data <= 32'hBE274336;	14'h1C31: data <= 32'hBE76F32A;	14'h1C32: data <= 32'hBEC6A31E;	14'h1C33: data <= 32'hBF165312;	14'h1C34: data <= 32'hBF660306;	14'h1C35: data <= 32'hBFB5B2FA;	14'h1C36: data <= 32'hC00562ED;	14'h1C37: data <= 32'hC05512E1;	14'h1C38: data <= 32'hC0A4C2D5;	14'h1C39: data <= 32'hC0F472C9;	14'h1C3A: data <= 32'hC14422BD;	14'h1C3B: data <= 32'hC193D2B1;	14'h1C3C: data <= 32'hC1E382A5;	14'h1C3D: data <= 32'hC2310263;	14'h1C3E: data <= 32'hC266BFD6;	14'h1C3F: data <= 32'hC29C7D49;	14'h1C40: data <= 32'hC2D23ABC;	14'h1C41: data <= 32'hC307F82F;	14'h1C42: data <= 32'hC33DB5A3;	14'h1C43: data <= 32'hC3737316;	14'h1C44: data <= 32'hC3A93089;	14'h1C45: data <= 32'hC3DEEDFC;	14'h1C46: data <= 32'hC414AB6F;	14'h1C47: data <= 32'hC44A68E2;	14'h1C48: data <= 32'hC4802656;	14'h1C49: data <= 32'hC4B5E3C9;	14'h1C4A: data <= 32'hC4EBA13C;	14'h1C4B: data <= 32'hC5215EAF;	14'h1C4C: data <= 32'hC5571C22;	14'h1C4D: data <= 32'hC58CD995;	14'h1C4E: data <= 32'hC5C29708;	14'h1C4F: data <= 32'hC5F8547C;	14'h1C50: data <= 32'hC62E11EF;	14'h1C51: data <= 32'hC663CF62;	14'h1C52: data <= 32'hC6998CD5;	14'h1C53: data <= 32'hC6CF4A48;	14'h1C54: data <= 32'hC70507BB;	14'h1C55: data <= 32'hC73AC52F;	14'h1C56: data <= 32'hC77082A2;	14'h1C57: data <= 32'hC7A64015;	14'h1C58: data <= 32'hC7DBFD88;	14'h1C59: data <= 32'hC811BAFB;	14'h1C5A: data <= 32'hC847786E;	14'h1C5B: data <= 32'hC87D35E1;	14'h1C5C: data <= 32'hC8B2F355;	14'h1C5D: data <= 32'hC8E8B0C8;	14'h1C5E: data <= 32'hC91E6E3B;	14'h1C5F: data <= 32'hC9542BAE;	14'h1C60: data <= 32'hC989E921;	14'h1C61: data <= 32'hC9BFA694;	14'h1C62: data <= 32'hC9F498CD;	14'h1C63: data <= 32'hCA297DFF;	14'h1C64: data <= 32'hCA5E6331;	14'h1C65: data <= 32'hCA934863;	14'h1C66: data <= 32'hCAC82D95;	14'h1C67: data <= 32'hCAFD12C7;	14'h1C68: data <= 32'hCB31F7F9;	14'h1C69: data <= 32'hCB66DD2B;	14'h1C6A: data <= 32'hCB9BC25D;	14'h1C6B: data <= 32'hCBD0A78F;	14'h1C6C: data <= 32'hCC058CC1;	14'h1C6D: data <= 32'hCC3A71F3;	14'h1C6E: data <= 32'hCC6F5725;	14'h1C6F: data <= 32'hCCA43C57;	14'h1C70: data <= 32'hCCD92188;	14'h1C71: data <= 32'hCD0E06BA;	14'h1C72: data <= 32'hCD42EBEC;	14'h1C73: data <= 32'hCD77D11E;	14'h1C74: data <= 32'hCDACB650;	14'h1C75: data <= 32'hCDE19B82;	14'h1C76: data <= 32'hCE1680B4;	14'h1C77: data <= 32'hCE4B65E6;	14'h1C78: data <= 32'hCE804B18;	14'h1C79: data <= 32'hCEB5304A;	14'h1C7A: data <= 32'hCEEA157C;	14'h1C7B: data <= 32'hCF1EFAAE;	14'h1C7C: data <= 32'hCF53DFE0;	14'h1C7D: data <= 32'hCF88C512;	14'h1C7E: data <= 32'hCFBDAA44;	14'h1C7F: data <= 32'hCFF28F75;	14'h1C80: data <= 32'hD02774A7;	14'h1C81: data <= 32'hD05C59D9;	14'h1C82: data <= 32'hD0913F0B;	14'h1C83: data <= 32'hD0C6243D;	14'h1C84: data <= 32'hD0FB096F;	14'h1C85: data <= 32'hD12FEEA1;	14'h1C86: data <= 32'hD167123C;	14'h1C87: data <= 32'hD19EC9CC;	14'h1C88: data <= 32'hD1D6815B;	14'h1C89: data <= 32'hD20E38EB;	14'h1C8A: data <= 32'hD245F07A;	14'h1C8B: data <= 32'hD27DA80A;	14'h1C8C: data <= 32'hD2B55F99;	14'h1C8D: data <= 32'hD2ED1729;	14'h1C8E: data <= 32'hD324CEB8;	14'h1C8F: data <= 32'hD35C8648;	14'h1C90: data <= 32'hD3943DD7;	14'h1C91: data <= 32'hD3CBF567;	14'h1C92: data <= 32'hD403ACF6;	14'h1C93: data <= 32'hD43B6486;	14'h1C94: data <= 32'hD4731C15;	14'h1C95: data <= 32'hD4AAD3A5;	14'h1C96: data <= 32'hD4E28B34;	14'h1C97: data <= 32'hD51A42C4;	14'h1C98: data <= 32'hD551FA53;	14'h1C99: data <= 32'hD589B1E3;	14'h1C9A: data <= 32'hD5C16972;	14'h1C9B: data <= 32'hD5F92102;	14'h1C9C: data <= 32'hD630D892;	14'h1C9D: data <= 32'hD6689021;	14'h1C9E: data <= 32'hD6A047B1;	14'h1C9F: data <= 32'hD6D7FF40;	14'h1CA0: data <= 32'hD70FB6D0;	14'h1CA1: data <= 32'hD7476E5F;	14'h1CA2: data <= 32'hD77F25EF;	14'h1CA3: data <= 32'hD7B6DD7E;	14'h1CA4: data <= 32'hD7EE950E;	14'h1CA5: data <= 32'hD8264C9D;	14'h1CA6: data <= 32'hD85E042D;	14'h1CA7: data <= 32'hD895BBBC;	14'h1CA8: data <= 32'hD8CD734C;	14'h1CA9: data <= 32'hD9052ADB;	14'h1CAA: data <= 32'hD93BA699;	14'h1CAB: data <= 32'hD97178BD;	14'h1CAC: data <= 32'hD9A74AE0;	14'h1CAD: data <= 32'hD9DD1D03;	14'h1CAE: data <= 32'hDA12EF27;	14'h1CAF: data <= 32'hDA48C14A;	14'h1CB0: data <= 32'hDA7E936D;	14'h1CB1: data <= 32'hDAB46591;	14'h1CB2: data <= 32'hDAEA37B4;	14'h1CB3: data <= 32'hDB2009D7;	14'h1CB4: data <= 32'hDB55DBFB;	14'h1CB5: data <= 32'hDB8BAE1E;	14'h1CB6: data <= 32'hDBC18041;	14'h1CB7: data <= 32'hDBF75265;	14'h1CB8: data <= 32'hDC2D2488;	14'h1CB9: data <= 32'hDC62F6AB;	14'h1CBA: data <= 32'hDC98C8CF;	14'h1CBB: data <= 32'hDCCE9AF2;	14'h1CBC: data <= 32'hDD046D15;	14'h1CBD: data <= 32'hDD3A3F39;	14'h1CBE: data <= 32'hDD70115C;	14'h1CBF: data <= 32'hDDA5E37F;	14'h1CC0: data <= 32'hDDDBB5A3;	14'h1CC1: data <= 32'hDE1187C6;	14'h1CC2: data <= 32'hDE4759E9;	14'h1CC3: data <= 32'hDE7D2C0D;	14'h1CC4: data <= 32'hDEB2FE30;	14'h1CC5: data <= 32'hDEE8D053;	14'h1CC6: data <= 32'hDF1EA277;	14'h1CC7: data <= 32'hDF54749A;	14'h1CC8: data <= 32'hDF8A46BD;	14'h1CC9: data <= 32'hDFC018E1;	14'h1CCA: data <= 32'hDFF5EB04;	14'h1CCB: data <= 32'hE02BBD27;	14'h1CCC: data <= 32'hE0618F4B;	14'h1CCD: data <= 32'hE097616E;	14'h1CCE: data <= 32'hE0C5673F;	14'h1CCF: data <= 32'hE0EBD045;	14'h1CD0: data <= 32'hE112394C;	14'h1CD1: data <= 32'hE138A252;	14'h1CD2: data <= 32'hE15F0B59;	14'h1CD3: data <= 32'hE185745F;	14'h1CD4: data <= 32'hE1ABDD66;	14'h1CD5: data <= 32'hE1D2466C;	14'h1CD6: data <= 32'hE1F8AF73;	14'h1CD7: data <= 32'hE21F1879;	14'h1CD8: data <= 32'hE2458180;	14'h1CD9: data <= 32'hE26BEA86;	14'h1CDA: data <= 32'hE292538C;	14'h1CDB: data <= 32'hE2B8BC93;	14'h1CDC: data <= 32'hE2DF2599;	14'h1CDD: data <= 32'hE3058EA0;	14'h1CDE: data <= 32'hE32BF7A6;	14'h1CDF: data <= 32'hE35260AD;	14'h1CE0: data <= 32'hE378C9B3;	14'h1CE1: data <= 32'hE39F32BA;	14'h1CE2: data <= 32'hE3C59BC0;	14'h1CE3: data <= 32'hE3EC04C7;	14'h1CE4: data <= 32'hE4126DCD;	14'h1CE5: data <= 32'hE438D6D4;	14'h1CE6: data <= 32'hE45F3FDA;	14'h1CE7: data <= 32'hE485A8E0;	14'h1CE8: data <= 32'hE4AC11E7;	14'h1CE9: data <= 32'hE4D27AED;	14'h1CEA: data <= 32'hE4F8E3F4;	14'h1CEB: data <= 32'hE51F4CFA;	14'h1CEC: data <= 32'hE545B601;	14'h1CED: data <= 32'hE56C1F07;	14'h1CEE: data <= 32'hE592880E;	14'h1CEF: data <= 32'hE5B8F114;	14'h1CF0: data <= 32'hE5DF5A1B;	14'h1CF1: data <= 32'hE605C321;	14'h1CF2: data <= 32'hE6280F4F;	14'h1CF3: data <= 32'hE6431778;	14'h1CF4: data <= 32'hE65E1FA0;	14'h1CF5: data <= 32'hE67927C8;	14'h1CF6: data <= 32'hE6942FF0;	14'h1CF7: data <= 32'hE6AF3818;	14'h1CF8: data <= 32'hE6CA4040;	14'h1CF9: data <= 32'hE6E54868;	14'h1CFA: data <= 32'hE7005090;	14'h1CFB: data <= 32'hE71B58B8;	14'h1CFC: data <= 32'hE73660E0;	14'h1CFD: data <= 32'hE7516909;	14'h1CFE: data <= 32'hE76C7131;	14'h1CFF: data <= 32'hE7877959;	14'h1D00: data <= 32'hE7A28181;	14'h1D01: data <= 32'hE7BD89A9;	14'h1D02: data <= 32'hE7D891D1;	14'h1D03: data <= 32'hE7F399F9;	14'h1D04: data <= 32'hE80EA221;	14'h1D05: data <= 32'hE829AA49;	14'h1D06: data <= 32'hE844B272;	14'h1D07: data <= 32'hE85FBA9A;	14'h1D08: data <= 32'hE87AC2C2;	14'h1D09: data <= 32'hE895CAEA;	14'h1D0A: data <= 32'hE8B0D312;	14'h1D0B: data <= 32'hE8CBDB3A;	14'h1D0C: data <= 32'hE8E6E362;	14'h1D0D: data <= 32'hE901EB8A;	14'h1D0E: data <= 32'hE91CF3B2;	14'h1D0F: data <= 32'hE937FBDB;	14'h1D10: data <= 32'hE9530403;	14'h1D11: data <= 32'hE96E0C2B;	14'h1D12: data <= 32'hE9891453;	14'h1D13: data <= 32'hE9A41C7B;	14'h1D14: data <= 32'hE9BF24A3;	14'h1D15: data <= 32'hE9DA2CCB;	14'h1D16: data <= 32'hE9F2AF3E;	14'h1D17: data <= 32'hEA0215F8;	14'h1D18: data <= 32'hEA117CB3;	14'h1D19: data <= 32'hEA20E36D;	14'h1D1A: data <= 32'hEA304A27;	14'h1D1B: data <= 32'hEA3FB0E2;	14'h1D1C: data <= 32'hEA4F179C;	14'h1D1D: data <= 32'hEA5E7E56;	14'h1D1E: data <= 32'hEA6DE511;	14'h1D1F: data <= 32'hEA7D4BCB;	14'h1D20: data <= 32'hEA8CB285;	14'h1D21: data <= 32'hEA9C1940;	14'h1D22: data <= 32'hEAAB7FFA;	14'h1D23: data <= 32'hEABAE6B4;	14'h1D24: data <= 32'hEACA4D6F;	14'h1D25: data <= 32'hEAD9B429;	14'h1D26: data <= 32'hEAE91AE3;	14'h1D27: data <= 32'hEAF8819E;	14'h1D28: data <= 32'hEB07E858;	14'h1D29: data <= 32'hEB174F12;	14'h1D2A: data <= 32'hEB26B5CD;	14'h1D2B: data <= 32'hEB361C87;	14'h1D2C: data <= 32'hEB458341;	14'h1D2D: data <= 32'hEB54E9FC;	14'h1D2E: data <= 32'hEB6450B6;	14'h1D2F: data <= 32'hEB73B770;	14'h1D30: data <= 32'hEB831E2B;	14'h1D31: data <= 32'hEB9284E5;	14'h1D32: data <= 32'hEBA1EB9F;	14'h1D33: data <= 32'hEBB15259;	14'h1D34: data <= 32'hEBC0B914;	14'h1D35: data <= 32'hEBD01FCE;	14'h1D36: data <= 32'hEBDF8688;	14'h1D37: data <= 32'hEBEEED43;	14'h1D38: data <= 32'hEBFE53FD;	14'h1D39: data <= 32'hEC0DBAB7;	14'h1D3A: data <= 32'hEC1C0FA4;	14'h1D3B: data <= 32'hEC1CAAC7;	14'h1D3C: data <= 32'hEC1D45E9;	14'h1D3D: data <= 32'hEC1DE10B;	14'h1D3E: data <= 32'hEC1E7C2D;	14'h1D3F: data <= 32'hEC1F174F;	14'h1D40: data <= 32'hEC1FB271;	14'h1D41: data <= 32'hEC204D93;	14'h1D42: data <= 32'hEC20E8B6;	14'h1D43: data <= 32'hEC2183D8;	14'h1D44: data <= 32'hEC221EFA;	14'h1D45: data <= 32'hEC22BA1C;	14'h1D46: data <= 32'hEC23553E;	14'h1D47: data <= 32'hEC23F060;	14'h1D48: data <= 32'hEC248B82;	14'h1D49: data <= 32'hEC2526A5;	14'h1D4A: data <= 32'hEC25C1C7;	14'h1D4B: data <= 32'hEC265CE9;	14'h1D4C: data <= 32'hEC26F80B;	14'h1D4D: data <= 32'hEC27932D;	14'h1D4E: data <= 32'hEC282E4F;	14'h1D4F: data <= 32'hEC28C971;	14'h1D50: data <= 32'hEC296494;	14'h1D51: data <= 32'hEC29FFB6;	14'h1D52: data <= 32'hEC2A9AD8;	14'h1D53: data <= 32'hEC2B35FA;	14'h1D54: data <= 32'hEC2BD11C;	14'h1D55: data <= 32'hEC2C6C3E;	14'h1D56: data <= 32'hEC2D0760;	14'h1D57: data <= 32'hEC2DA283;	14'h1D58: data <= 32'hEC2E3DA5;	14'h1D59: data <= 32'hEC2ED8C7;	14'h1D5A: data <= 32'hEC2F73E9;	14'h1D5B: data <= 32'hEC300F0B;	14'h1D5C: data <= 32'hEC30AA2D;	14'h1D5D: data <= 32'hEC31454F;	14'h1D5E: data <= 32'hEC31E072;	14'h1D5F: data <= 32'hEC2DFDFA;	14'h1D60: data <= 32'hEC29C1ED;	14'h1D61: data <= 32'hEC2585E1;	14'h1D62: data <= 32'hEC2149D5;	14'h1D63: data <= 32'hEC1D0DC9;	14'h1D64: data <= 32'hEC18D1BD;	14'h1D65: data <= 32'hEC1495B0;	14'h1D66: data <= 32'hEC1059A4;	14'h1D67: data <= 32'hEC0C1D98;	14'h1D68: data <= 32'hEC07E18C;	14'h1D69: data <= 32'hEC03A57F;	14'h1D6A: data <= 32'hEBFF6973;	14'h1D6B: data <= 32'hEBFB2D67;	14'h1D6C: data <= 32'hEBF6F15B;	14'h1D6D: data <= 32'hEBF2B54F;	14'h1D6E: data <= 32'hEBEE7942;	14'h1D6F: data <= 32'hEBEA3D36;	14'h1D70: data <= 32'hEBE6012A;	14'h1D71: data <= 32'hEBE1C51E;	14'h1D72: data <= 32'hEBDD8911;	14'h1D73: data <= 32'hEBD94D05;	14'h1D74: data <= 32'hEBD510F9;	14'h1D75: data <= 32'hEBD0D4ED;	14'h1D76: data <= 32'hEBCC98E0;	14'h1D77: data <= 32'hEBC85CD4;	14'h1D78: data <= 32'hEBC420C8;	14'h1D79: data <= 32'hEBBFE4BC;	14'h1D7A: data <= 32'hEBBBA8B0;	14'h1D7B: data <= 32'hEBB76CA3;	14'h1D7C: data <= 32'hEBB33097;	14'h1D7D: data <= 32'hEBAEF48B;	14'h1D7E: data <= 32'hEBAAB87F;	14'h1D7F: data <= 32'hEBA67C72;	14'h1D80: data <= 32'hEBA24066;	14'h1D81: data <= 32'hEB9E045A;	14'h1D82: data <= 32'hEB99C84E;	14'h1D83: data <= 32'hEB9D59D3;	14'h1D84: data <= 32'hEBA31485;	14'h1D85: data <= 32'hEBA8CF37;	14'h1D86: data <= 32'hEBAE89E9;	14'h1D87: data <= 32'hEBB4449B;	14'h1D88: data <= 32'hEBB9FF4D;	14'h1D89: data <= 32'hEBBFB9FF;	14'h1D8A: data <= 32'hEBC574B1;	14'h1D8B: data <= 32'hEBCB2F63;	14'h1D8C: data <= 32'hEBD0EA15;	14'h1D8D: data <= 32'hEBD6A4C7;	14'h1D8E: data <= 32'hEBDC5F79;	14'h1D8F: data <= 32'hEBE21A2B;	14'h1D90: data <= 32'hEBE7D4DD;	14'h1D91: data <= 32'hEBED8F8F;	14'h1D92: data <= 32'hEBF34A41;	14'h1D93: data <= 32'hEBF904F3;	14'h1D94: data <= 32'hEBFEBFA5;	14'h1D95: data <= 32'hEC047A57;	14'h1D96: data <= 32'hEC0A3509;	14'h1D97: data <= 32'hEC0FEFBB;	14'h1D98: data <= 32'hEC15AA6D;	14'h1D99: data <= 32'hEC1B651F;	14'h1D9A: data <= 32'hEC211FD0;	14'h1D9B: data <= 32'hEC26DA82;	14'h1D9C: data <= 32'hEC2C9534;	14'h1D9D: data <= 32'hEC324FE6;	14'h1D9E: data <= 32'hEC380A98;	14'h1D9F: data <= 32'hEC3DC54A;	14'h1DA0: data <= 32'hEC437FFC;	14'h1DA1: data <= 32'hEC493AAE;	14'h1DA2: data <= 32'hEC4EF560;	14'h1DA3: data <= 32'hEC54B012;	14'h1DA4: data <= 32'hEC5A6AC4;	14'h1DA5: data <= 32'hEC602576;	14'h1DA6: data <= 32'hEC65E028;	14'h1DA7: data <= 32'hEC7000F8;	14'h1DA8: data <= 32'hEC7C9F34;	14'h1DA9: data <= 32'hEC893D70;	14'h1DAA: data <= 32'hEC95DBAC;	14'h1DAB: data <= 32'hECA279E8;	14'h1DAC: data <= 32'hECAF1824;	14'h1DAD: data <= 32'hECBBB660;	14'h1DAE: data <= 32'hECC8549C;	14'h1DAF: data <= 32'hECD4F2D8;	14'h1DB0: data <= 32'hECE19114;	14'h1DB1: data <= 32'hECEE2F51;	14'h1DB2: data <= 32'hECFACD8D;	14'h1DB3: data <= 32'hED076BC9;	14'h1DB4: data <= 32'hED140A05;	14'h1DB5: data <= 32'hED20A841;	14'h1DB6: data <= 32'hED2D467D;	14'h1DB7: data <= 32'hED39E4B9;	14'h1DB8: data <= 32'hED4682F5;	14'h1DB9: data <= 32'hED532131;	14'h1DBA: data <= 32'hED5FBF6D;	14'h1DBB: data <= 32'hED6C5DA9;	14'h1DBC: data <= 32'hED78FBE6;	14'h1DBD: data <= 32'hED859A22;	14'h1DBE: data <= 32'hED92385E;	14'h1DBF: data <= 32'hED9ED69A;	14'h1DC0: data <= 32'hEDAB74D6;	14'h1DC1: data <= 32'hEDB81312;	14'h1DC2: data <= 32'hEDC4B14E;	14'h1DC3: data <= 32'hEDD14F8A;	14'h1DC4: data <= 32'hEDDDEDC6;	14'h1DC5: data <= 32'hEDEA8C02;	14'h1DC6: data <= 32'hEDF72A3F;	14'h1DC7: data <= 32'hEE03C87B;	14'h1DC8: data <= 32'hEE1066B7;	14'h1DC9: data <= 32'hEE1D04F3;	14'h1DCA: data <= 32'hEE29A32F;	14'h1DCB: data <= 32'hEE361660;	14'h1DCC: data <= 32'hEE425D7A;	14'h1DCD: data <= 32'hEE4EA494;	14'h1DCE: data <= 32'hEE5AEBAD;	14'h1DCF: data <= 32'hEE6732C7;	14'h1DD0: data <= 32'hEE7379E1;	14'h1DD1: data <= 32'hEE7FC0FB;	14'h1DD2: data <= 32'hEE8C0814;	14'h1DD3: data <= 32'hEE984F2E;	14'h1DD4: data <= 32'hEEA49648;	14'h1DD5: data <= 32'hEEB0DD62;	14'h1DD6: data <= 32'hEEBD247B;	14'h1DD7: data <= 32'hEEC96B95;	14'h1DD8: data <= 32'hEED5B2AF;	14'h1DD9: data <= 32'hEEE1F9C8;	14'h1DDA: data <= 32'hEEEE40E2;	14'h1DDB: data <= 32'hEEFA87FC;	14'h1DDC: data <= 32'hEF06CF16;	14'h1DDD: data <= 32'hEF13162F;	14'h1DDE: data <= 32'hEF1F5D49;	14'h1DDF: data <= 32'hEF2BA463;	14'h1DE0: data <= 32'hEF37EB7D;	14'h1DE1: data <= 32'hEF443296;	14'h1DE2: data <= 32'hEF5079B0;	14'h1DE3: data <= 32'hEF5CC0CA;	14'h1DE4: data <= 32'hEF6907E4;	14'h1DE5: data <= 32'hEF754EFD;	14'h1DE6: data <= 32'hEF819617;	14'h1DE7: data <= 32'hEF8DDD31;	14'h1DE8: data <= 32'hEF9A244A;	14'h1DE9: data <= 32'hEFA66B64;	14'h1DEA: data <= 32'hEFB2B27E;	14'h1DEB: data <= 32'hEFBEF998;	14'h1DEC: data <= 32'hEFCB40B1;	14'h1DED: data <= 32'hEFD787CB;	14'h1DEE: data <= 32'hEFE3CEE5;	14'h1DEF: data <= 32'hEFF0CDF1;	14'h1DF0: data <= 32'hEFFF2382;	14'h1DF1: data <= 32'hF00D7913;	14'h1DF2: data <= 32'hF01BCEA4;	14'h1DF3: data <= 32'hF02A2435;	14'h1DF4: data <= 32'hF03879C6;	14'h1DF5: data <= 32'hF046CF57;	14'h1DF6: data <= 32'hF05524E8;	14'h1DF7: data <= 32'hF0637A79;	14'h1DF8: data <= 32'hF071D00A;	14'h1DF9: data <= 32'hF080259B;	14'h1DFA: data <= 32'hF08E7B2C;	14'h1DFB: data <= 32'hF09CD0BD;	14'h1DFC: data <= 32'hF0AB264E;	14'h1DFD: data <= 32'hF0B97BDF;	14'h1DFE: data <= 32'hF0C7D171;	14'h1DFF: data <= 32'hF0D62702;	14'h1E00: data <= 32'hF0E47C93;	14'h1E01: data <= 32'hF0F2D224;	14'h1E02: data <= 32'hF10127B5;	14'h1E03: data <= 32'hF10F7D46;	14'h1E04: data <= 32'hF11DD2D7;	14'h1E05: data <= 32'hF12C2868;	14'h1E06: data <= 32'hF13A7DF9;	14'h1E07: data <= 32'hF148D38A;	14'h1E08: data <= 32'hF157291B;	14'h1E09: data <= 32'hF1657EAC;	14'h1E0A: data <= 32'hF173D43D;	14'h1E0B: data <= 32'hF18229CE;	14'h1E0C: data <= 32'hF1907F5F;	14'h1E0D: data <= 32'hF19ED4F0;	14'h1E0E: data <= 32'hF1AD2A81;	14'h1E0F: data <= 32'hF1BB8012;	14'h1E10: data <= 32'hF1C9D5A3;	14'h1E11: data <= 32'hF1D82B34;	14'h1E12: data <= 32'hF1E680C6;	14'h1E13: data <= 32'hF1F55033;	14'h1E14: data <= 32'hF205F8BB;	14'h1E15: data <= 32'hF216A143;	14'h1E16: data <= 32'hF22749CB;	14'h1E17: data <= 32'hF237F253;	14'h1E18: data <= 32'hF2489ADB;	14'h1E19: data <= 32'hF2594362;	14'h1E1A: data <= 32'hF269EBEA;	14'h1E1B: data <= 32'hF27A9472;	14'h1E1C: data <= 32'hF28B3CFA;	14'h1E1D: data <= 32'hF29BE582;	14'h1E1E: data <= 32'hF2AC8E0A;	14'h1E1F: data <= 32'hF2BD3692;	14'h1E20: data <= 32'hF2CDDF1A;	14'h1E21: data <= 32'hF2DE87A2;	14'h1E22: data <= 32'hF2EF302A;	14'h1E23: data <= 32'hF2FFD8B2;	14'h1E24: data <= 32'hF310813A;	14'h1E25: data <= 32'hF32129C2;	14'h1E26: data <= 32'hF331D24A;	14'h1E27: data <= 32'hF3427AD2;	14'h1E28: data <= 32'hF353235A;	14'h1E29: data <= 32'hF363CBE2;	14'h1E2A: data <= 32'hF3747469;	14'h1E2B: data <= 32'hF3851CF1;	14'h1E2C: data <= 32'hF395C579;	14'h1E2D: data <= 32'hF3A66E01;	14'h1E2E: data <= 32'hF3B71689;	14'h1E2F: data <= 32'hF3C7BF11;	14'h1E30: data <= 32'hF3D86799;	14'h1E31: data <= 32'hF3E91021;	14'h1E32: data <= 32'hF3F9B8A9;	14'h1E33: data <= 32'hF40A6131;	14'h1E34: data <= 32'hF41B09B9;	14'h1E35: data <= 32'hF42BB241;	14'h1E36: data <= 32'hF43C5AC9;	14'h1E37: data <= 32'hF44CACDD;	14'h1E38: data <= 32'hF457BA51;	14'h1E39: data <= 32'hF462C7C4;	14'h1E3A: data <= 32'hF46DD537;	14'h1E3B: data <= 32'hF478E2AB;	14'h1E3C: data <= 32'hF483F01E;	14'h1E3D: data <= 32'hF48EFD91;	14'h1E3E: data <= 32'hF49A0B05;	14'h1E3F: data <= 32'hF4A51878;	14'h1E40: data <= 32'hF4B025EB;	14'h1E41: data <= 32'hF4BB335F;	14'h1E42: data <= 32'hF4C640D2;	14'h1E43: data <= 32'hF4D14E45;	14'h1E44: data <= 32'hF4DC5BB8;	14'h1E45: data <= 32'hF4E7692C;	14'h1E46: data <= 32'hF4F2769F;	14'h1E47: data <= 32'hF4FD8412;	14'h1E48: data <= 32'hF5089186;	14'h1E49: data <= 32'hF5139EF9;	14'h1E4A: data <= 32'hF51EAC6C;	14'h1E4B: data <= 32'hF529B9E0;	14'h1E4C: data <= 32'hF534C753;	14'h1E4D: data <= 32'hF53FD4C6;	14'h1E4E: data <= 32'hF54AE23A;	14'h1E4F: data <= 32'hF555EFAD;	14'h1E50: data <= 32'hF560FD20;	14'h1E51: data <= 32'hF56C0A94;	14'h1E52: data <= 32'hF5771807;	14'h1E53: data <= 32'hF582257A;	14'h1E54: data <= 32'hF58D32ED;	14'h1E55: data <= 32'hF5984061;	14'h1E56: data <= 32'hF5A34DD4;	14'h1E57: data <= 32'hF5AE5B47;	14'h1E58: data <= 32'hF5B968BB;	14'h1E59: data <= 32'hF5C4762E;	14'h1E5A: data <= 32'hF5CF83A1;	14'h1E5B: data <= 32'hF5DA9115;	14'h1E5C: data <= 32'hF5E02A28;	14'h1E5D: data <= 32'hF5E5429E;	14'h1E5E: data <= 32'hF5EA5B15;	14'h1E5F: data <= 32'hF5EF738B;	14'h1E60: data <= 32'hF5F48C02;	14'h1E61: data <= 32'hF5F9A478;	14'h1E62: data <= 32'hF5FEBCEE;	14'h1E63: data <= 32'hF603D565;	14'h1E64: data <= 32'hF608EDDB;	14'h1E65: data <= 32'hF60E0651;	14'h1E66: data <= 32'hF6131EC8;	14'h1E67: data <= 32'hF618373E;	14'h1E68: data <= 32'hF61D4FB4;	14'h1E69: data <= 32'hF622682B;	14'h1E6A: data <= 32'hF62780A1;	14'h1E6B: data <= 32'hF62C9918;	14'h1E6C: data <= 32'hF631B18E;	14'h1E6D: data <= 32'hF636CA04;	14'h1E6E: data <= 32'hF63BE27B;	14'h1E6F: data <= 32'hF640FAF1;	14'h1E70: data <= 32'hF6461367;	14'h1E71: data <= 32'hF64B2BDE;	14'h1E72: data <= 32'hF6504454;	14'h1E73: data <= 32'hF6555CCA;	14'h1E74: data <= 32'hF65A7541;	14'h1E75: data <= 32'hF65F8DB7;	14'h1E76: data <= 32'hF664A62E;	14'h1E77: data <= 32'hF669BEA4;	14'h1E78: data <= 32'hF66ED71A;	14'h1E79: data <= 32'hF673EF91;	14'h1E7A: data <= 32'hF6790807;	14'h1E7B: data <= 32'hF67E207D;	14'h1E7C: data <= 32'hF68338F4;	14'h1E7D: data <= 32'hF688516A;	14'h1E7E: data <= 32'hF68D69E0;	14'h1E7F: data <= 32'hF6928257;	14'h1E80: data <= 32'hF695FFCE;	14'h1E81: data <= 32'hF6990342;	14'h1E82: data <= 32'hF69C06B5;	14'h1E83: data <= 32'hF69F0A29;	14'h1E84: data <= 32'hF6A20D9C;	14'h1E85: data <= 32'hF6A51110;	14'h1E86: data <= 32'hF6A81484;	14'h1E87: data <= 32'hF6AB17F7;	14'h1E88: data <= 32'hF6AE1B6B;	14'h1E89: data <= 32'hF6B11EDE;	14'h1E8A: data <= 32'hF6B42252;	14'h1E8B: data <= 32'hF6B725C6;	14'h1E8C: data <= 32'hF6BA2939;	14'h1E8D: data <= 32'hF6BD2CAD;	14'h1E8E: data <= 32'hF6C03020;	14'h1E8F: data <= 32'hF6C33394;	14'h1E90: data <= 32'hF6C63707;	14'h1E91: data <= 32'hF6C93A7B;	14'h1E92: data <= 32'hF6CC3DEF;	14'h1E93: data <= 32'hF6CF4162;	14'h1E94: data <= 32'hF6D244D6;	14'h1E95: data <= 32'hF6D54849;	14'h1E96: data <= 32'hF6D84BBD;	14'h1E97: data <= 32'hF6DB4F31;	14'h1E98: data <= 32'hF6DE52A4;	14'h1E99: data <= 32'hF6E15618;	14'h1E9A: data <= 32'hF6E4598B;	14'h1E9B: data <= 32'hF6E75CFF;	14'h1E9C: data <= 32'hF6EA6072;	14'h1E9D: data <= 32'hF6ED63E6;	14'h1E9E: data <= 32'hF6F0675A;	14'h1E9F: data <= 32'hF6F36ACD;	14'h1EA0: data <= 32'hF6F66E41;	14'h1EA1: data <= 32'hF6F971B4;	14'h1EA2: data <= 32'hF6FC7528;	14'h1EA3: data <= 32'hF6FF789C;	14'h1EA4: data <= 32'hF7011868;	14'h1EA5: data <= 32'hF701E42F;	14'h1EA6: data <= 32'hF702AFF5;	14'h1EA7: data <= 32'hF7037BBC;	14'h1EA8: data <= 32'hF7044782;	14'h1EA9: data <= 32'hF7051349;	14'h1EAA: data <= 32'hF705DF0F;	14'h1EAB: data <= 32'hF706AAD6;	14'h1EAC: data <= 32'hF707769C;	14'h1EAD: data <= 32'hF7084263;	14'h1EAE: data <= 32'hF7090E29;	14'h1EAF: data <= 32'hF709D9F0;	14'h1EB0: data <= 32'hF70AA5B6;	14'h1EB1: data <= 32'hF70B717D;	14'h1EB2: data <= 32'hF70C3D43;	14'h1EB3: data <= 32'hF70D090A;	14'h1EB4: data <= 32'hF70DD4D1;	14'h1EB5: data <= 32'hF70EA097;	14'h1EB6: data <= 32'hF70F6C5E;	14'h1EB7: data <= 32'hF7103824;	14'h1EB8: data <= 32'hF71103EB;	14'h1EB9: data <= 32'hF711CFB1;	14'h1EBA: data <= 32'hF7129B78;	14'h1EBB: data <= 32'hF713673E;	14'h1EBC: data <= 32'hF7143305;	14'h1EBD: data <= 32'hF714FECB;	14'h1EBE: data <= 32'hF715CA92;	14'h1EBF: data <= 32'hF7169658;	14'h1EC0: data <= 32'hF717621F;	14'h1EC1: data <= 32'hF7182DE5;	14'h1EC2: data <= 32'hF718F9AC;	14'h1EC3: data <= 32'hF719C572;	14'h1EC4: data <= 32'hF71A9139;	14'h1EC5: data <= 32'hF71B5CFF;	14'h1EC6: data <= 32'hF71C28C6;	14'h1EC7: data <= 32'hF71CF48C;	14'h1EC8: data <= 32'hF71E31FB;	14'h1EC9: data <= 32'hF71FE997;	14'h1ECA: data <= 32'hF721A133;	14'h1ECB: data <= 32'hF72358CE;	14'h1ECC: data <= 32'hF725106A;	14'h1ECD: data <= 32'hF726C806;	14'h1ECE: data <= 32'hF7287FA2;	14'h1ECF: data <= 32'hF72A373E;	14'h1ED0: data <= 32'hF72BEEDA;	14'h1ED1: data <= 32'hF72DA676;	14'h1ED2: data <= 32'hF72F5E12;	14'h1ED3: data <= 32'hF73115AE;	14'h1ED4: data <= 32'hF732CD4A;	14'h1ED5: data <= 32'hF73484E6;	14'h1ED6: data <= 32'hF7363C82;	14'h1ED7: data <= 32'hF737F41E;	14'h1ED8: data <= 32'hF739ABBA;	14'h1ED9: data <= 32'hF73B6356;	14'h1EDA: data <= 32'hF73D1AF2;	14'h1EDB: data <= 32'hF73ED28E;	14'h1EDC: data <= 32'hF7408A2A;	14'h1EDD: data <= 32'hF74241C6;	14'h1EDE: data <= 32'hF743F961;	14'h1EDF: data <= 32'hF745B0FD;	14'h1EE0: data <= 32'hF7476899;	14'h1EE1: data <= 32'hF7492035;	14'h1EE2: data <= 32'hF74AD7D1;	14'h1EE3: data <= 32'hF74C8F6D;	14'h1EE4: data <= 32'hF74E4709;	14'h1EE5: data <= 32'hF74FFEA5;	14'h1EE6: data <= 32'hF751B641;	14'h1EE7: data <= 32'hF7536DDD;	14'h1EE8: data <= 32'hF7552579;	14'h1EE9: data <= 32'hF756DD15;	14'h1EEA: data <= 32'hF75894B1;	14'h1EEB: data <= 32'hF75A4C4D;	14'h1EEC: data <= 32'hF75C2E11;	14'h1EED: data <= 32'hF75E62A3;	14'h1EEE: data <= 32'hF7609734;	14'h1EEF: data <= 32'hF762CBC6;	14'h1EF0: data <= 32'hF7650058;	14'h1EF1: data <= 32'hF76734EA;	14'h1EF2: data <= 32'hF769697C;	14'h1EF3: data <= 32'hF76B9E0E;	14'h1EF4: data <= 32'hF76DD2A0;	14'h1EF5: data <= 32'hF7700732;	14'h1EF6: data <= 32'hF7723BC4;	14'h1EF7: data <= 32'hF7747056;	14'h1EF8: data <= 32'hF776A4E8;	14'h1EF9: data <= 32'hF778D97A;	14'h1EFA: data <= 32'hF77B0E0B;	14'h1EFB: data <= 32'hF77D429D;	14'h1EFC: data <= 32'hF77F772F;	14'h1EFD: data <= 32'hF781ABC1;	14'h1EFE: data <= 32'hF783E053;	14'h1EFF: data <= 32'hF78614E5;	14'h1F00: data <= 32'hF7884977;	14'h1F01: data <= 32'hF78A7E09;	14'h1F02: data <= 32'hF78CB29B;	14'h1F03: data <= 32'hF78EE72D;	14'h1F04: data <= 32'hF7911BBF;	14'h1F05: data <= 32'hF7935051;	14'h1F06: data <= 32'hF79584E2;	14'h1F07: data <= 32'hF797B974;	14'h1F08: data <= 32'hF799EE06;	14'h1F09: data <= 32'hF79C2298;	14'h1F0A: data <= 32'hF79E572A;	14'h1F0B: data <= 32'hF7A08BBC;	14'h1F0C: data <= 32'hF7A2C04E;	14'h1F0D: data <= 32'hF7A4F4E0;	14'h1F0E: data <= 32'hF7A72972;	14'h1F0F: data <= 32'hF7A95E04;	14'h1F10: data <= 32'hF7AB1572;	14'h1F11: data <= 32'hF7AAC0DD;	14'h1F12: data <= 32'hF7AA6C48;	14'h1F13: data <= 32'hF7AA17B3;	14'h1F14: data <= 32'hF7A9C31E;	14'h1F15: data <= 32'hF7A96E88;	14'h1F16: data <= 32'hF7A919F3;	14'h1F17: data <= 32'hF7A8C55E;	14'h1F18: data <= 32'hF7A870C9;	14'h1F19: data <= 32'hF7A81C34;	14'h1F1A: data <= 32'hF7A7C79E;	14'h1F1B: data <= 32'hF7A77309;	14'h1F1C: data <= 32'hF7A71E74;	14'h1F1D: data <= 32'hF7A6C9DF;	14'h1F1E: data <= 32'hF7A6754A;	14'h1F1F: data <= 32'hF7A620B4;	14'h1F20: data <= 32'hF7A5CC1F;	14'h1F21: data <= 32'hF7A5778A;	14'h1F22: data <= 32'hF7A522F5;	14'h1F23: data <= 32'hF7A4CE5F;	14'h1F24: data <= 32'hF7A479CA;	14'h1F25: data <= 32'hF7A42535;	14'h1F26: data <= 32'hF7A3D0A0;	14'h1F27: data <= 32'hF7A37C0B;	14'h1F28: data <= 32'hF7A32775;	14'h1F29: data <= 32'hF7A2D2E0;	14'h1F2A: data <= 32'hF7A27E4B;	14'h1F2B: data <= 32'hF7A229B6;	14'h1F2C: data <= 32'hF7A1D521;	14'h1F2D: data <= 32'hF7A1808B;	14'h1F2E: data <= 32'hF7A12BF6;	14'h1F2F: data <= 32'hF7A0D761;	14'h1F30: data <= 32'hF7A082CC;	14'h1F31: data <= 32'hF7A02E37;	14'h1F32: data <= 32'hF79FD9A1;	14'h1F33: data <= 32'hF79F850C;	14'h1F34: data <= 32'hF79F27FA;	14'h1F35: data <= 32'hF79E234C;	14'h1F36: data <= 32'hF79D1E9D;	14'h1F37: data <= 32'hF79C19EF;	14'h1F38: data <= 32'hF79B1540;	14'h1F39: data <= 32'hF79A1092;	14'h1F3A: data <= 32'hF7990BE3;	14'h1F3B: data <= 32'hF7980735;	14'h1F3C: data <= 32'hF7970286;	14'h1F3D: data <= 32'hF795FDD8;	14'h1F3E: data <= 32'hF794F929;	14'h1F3F: data <= 32'hF793F47B;	14'h1F40: data <= 32'hF792EFCC;	14'h1F41: data <= 32'hF791EB1E;	14'h1F42: data <= 32'hF790E66F;	14'h1F43: data <= 32'hF78FE1C1;	14'h1F44: data <= 32'hF78EDD12;	14'h1F45: data <= 32'hF78DD864;	14'h1F46: data <= 32'hF78CD3B5;	14'h1F47: data <= 32'hF78BCF07;	14'h1F48: data <= 32'hF78ACA58;	14'h1F49: data <= 32'hF789C5AA;	14'h1F4A: data <= 32'hF788C0FB;	14'h1F4B: data <= 32'hF787BC4C;	14'h1F4C: data <= 32'hF786B79E;	14'h1F4D: data <= 32'hF785B2EF;	14'h1F4E: data <= 32'hF784AE41;	14'h1F4F: data <= 32'hF783A992;	14'h1F50: data <= 32'hF782A4E4;	14'h1F51: data <= 32'hF781A035;	14'h1F52: data <= 32'hF7809B87;	14'h1F53: data <= 32'hF77F96D8;	14'h1F54: data <= 32'hF77E922A;	14'h1F55: data <= 32'hF77D8D7B;	14'h1F56: data <= 32'hF77C88CD;	14'h1F57: data <= 32'hF77B841E;	14'h1F58: data <= 32'hF77A7F70;	14'h1F59: data <= 32'hF774D10A;	14'h1F5A: data <= 32'hF76EA34F;	14'h1F5B: data <= 32'hF7687595;	14'h1F5C: data <= 32'hF76247DB;	14'h1F5D: data <= 32'hF75C1A20;	14'h1F5E: data <= 32'hF755EC66;	14'h1F5F: data <= 32'hF74FBEAC;	14'h1F60: data <= 32'hF74990F1;	14'h1F61: data <= 32'hF7436337;	14'h1F62: data <= 32'hF73D357D;	14'h1F63: data <= 32'hF73707C2;	14'h1F64: data <= 32'hF730DA08;	14'h1F65: data <= 32'hF72AAC4D;	14'h1F66: data <= 32'hF7247E93;	14'h1F67: data <= 32'hF71E50D9;	14'h1F68: data <= 32'hF718231E;	14'h1F69: data <= 32'hF711F564;	14'h1F6A: data <= 32'hF70BC7AA;	14'h1F6B: data <= 32'hF70599EF;	14'h1F6C: data <= 32'hF6FF6C35;	14'h1F6D: data <= 32'hF6F93E7B;	14'h1F6E: data <= 32'hF6F310C0;	14'h1F6F: data <= 32'hF6ECE306;	14'h1F70: data <= 32'hF6E6B54B;	14'h1F71: data <= 32'hF6E08791;	14'h1F72: data <= 32'hF6DA59D7;	14'h1F73: data <= 32'hF6D42C1C;	14'h1F74: data <= 32'hF6CDFE62;	14'h1F75: data <= 32'hF6C7D0A8;	14'h1F76: data <= 32'hF6C1A2ED;	14'h1F77: data <= 32'hF6BB7533;	14'h1F78: data <= 32'hF6B54779;	14'h1F79: data <= 32'hF6AF19BE;	14'h1F7A: data <= 32'hF6A8EC04;	14'h1F7B: data <= 32'hF6A2BE4A;	14'h1F7C: data <= 32'hF69C908F;	14'h1F7D: data <= 32'hF6912094;	14'h1F7E: data <= 32'hF6840538;	14'h1F7F: data <= 32'hF676E9DB;	14'h1F80: data <= 32'hF669CE7E;	14'h1F81: data <= 32'hF65CB322;	14'h1F82: data <= 32'hF64F97C5;	14'h1F83: data <= 32'hF6427C68;	14'h1F84: data <= 32'hF635610C;	14'h1F85: data <= 32'hF62845AF;	14'h1F86: data <= 32'hF61B2A52;	14'h1F87: data <= 32'hF60E0EF6;	14'h1F88: data <= 32'hF600F399;	14'h1F89: data <= 32'hF5F3D83C;	14'h1F8A: data <= 32'hF5E6BCE0;	14'h1F8B: data <= 32'hF5D9A183;	14'h1F8C: data <= 32'hF5CC8627;	14'h1F8D: data <= 32'hF5BF6ACA;	14'h1F8E: data <= 32'hF5B24F6D;	14'h1F8F: data <= 32'hF5A53411;	14'h1F90: data <= 32'hF59818B4;	14'h1F91: data <= 32'hF58AFD57;	14'h1F92: data <= 32'hF57DE1FB;	14'h1F93: data <= 32'hF570C69E;	14'h1F94: data <= 32'hF563AB41;	14'h1F95: data <= 32'hF5568FE5;	14'h1F96: data <= 32'hF5497488;	14'h1F97: data <= 32'hF53C592B;	14'h1F98: data <= 32'hF52F3DCF;	14'h1F99: data <= 32'hF5222272;	14'h1F9A: data <= 32'hF5150716;	14'h1F9B: data <= 32'hF507EBB9;	14'h1F9C: data <= 32'hF4FAD05C;	14'h1F9D: data <= 32'hF4EDB500;	14'h1F9E: data <= 32'hF4E099A3;	14'h1F9F: data <= 32'hF4D37E46;	14'h1FA0: data <= 32'hF4C662EA;	14'h1FA1: data <= 32'hF4B687FF;	14'h1FA2: data <= 32'hF4A4F3A1;	14'h1FA3: data <= 32'hF4935F44;	14'h1FA4: data <= 32'hF481CAE6;	14'h1FA5: data <= 32'hF4703689;	14'h1FA6: data <= 32'hF45EA22C;	14'h1FA7: data <= 32'hF44D0DCE;	14'h1FA8: data <= 32'hF43B7971;	14'h1FA9: data <= 32'hF429E514;	14'h1FAA: data <= 32'hF41850B6;	14'h1FAB: data <= 32'hF406BC59;	14'h1FAC: data <= 32'hF3F527FB;	14'h1FAD: data <= 32'hF3E3939E;	14'h1FAE: data <= 32'hF3D1FF41;	14'h1FAF: data <= 32'hF3C06AE3;	14'h1FB0: data <= 32'hF3AED686;	14'h1FB1: data <= 32'hF39D4228;	14'h1FB2: data <= 32'hF38BADCB;	14'h1FB3: data <= 32'hF37A196E;	14'h1FB4: data <= 32'hF3688510;	14'h1FB5: data <= 32'hF356F0B3;	14'h1FB6: data <= 32'hF3455C55;	14'h1FB7: data <= 32'hF333C7F8;	14'h1FB8: data <= 32'hF322339B;	14'h1FB9: data <= 32'hF3109F3D;	14'h1FBA: data <= 32'hF2FF0AE0;	14'h1FBB: data <= 32'hF2ED7682;	14'h1FBC: data <= 32'hF2DBE225;	14'h1FBD: data <= 32'hF2CA4DC8;	14'h1FBE: data <= 32'hF2B8B96A;	14'h1FBF: data <= 32'hF2A7250D;	14'h1FC0: data <= 32'hF29590AF;	14'h1FC1: data <= 32'hF283FC52;	14'h1FC2: data <= 32'hF27267F5;	14'h1FC3: data <= 32'hF260D397;	14'h1FC4: data <= 32'hF24F3F3A;	14'h1FC5: data <= 32'hF23CD87E;	14'h1FC6: data <= 32'hF229846C;	14'h1FC7: data <= 32'hF2163059;	14'h1FC8: data <= 32'hF202DC47;	14'h1FC9: data <= 32'hF1EF8835;	14'h1FCA: data <= 32'hF1DC3422;	14'h1FCB: data <= 32'hF1C8E010;	14'h1FCC: data <= 32'hF1B58BFE;	14'h1FCD: data <= 32'hF1A237EB;	14'h1FCE: data <= 32'hF18EE3D9;	14'h1FCF: data <= 32'hF17B8FC7;	14'h1FD0: data <= 32'hF1683BB4;	14'h1FD1: data <= 32'hF154E7A2;	14'h1FD2: data <= 32'hF1419390;	14'h1FD3: data <= 32'hF12E3F7D;	14'h1FD4: data <= 32'hF11AEB6B;	14'h1FD5: data <= 32'hF1079758;	14'h1FD6: data <= 32'hF0F44346;	14'h1FD7: data <= 32'hF0E0EF34;	14'h1FD8: data <= 32'hF0CD9B21;	14'h1FD9: data <= 32'hF0BA470F;	14'h1FDA: data <= 32'hF0A6F2FD;	14'h1FDB: data <= 32'hF0939EEA;	14'h1FDC: data <= 32'hF0804AD8;	14'h1FDD: data <= 32'hF06CF6C6;	14'h1FDE: data <= 32'hF059A2B3;	14'h1FDF: data <= 32'hF0464EA1;	14'h1FE0: data <= 32'hF032FA8F;	14'h1FE1: data <= 32'hF01FA67C;	14'h1FE2: data <= 32'hF00C526A;	14'h1FE3: data <= 32'hEFF8FE58;	14'h1FE4: data <= 32'hEFE5AA45;	14'h1FE5: data <= 32'hEFD25633;	14'h1FE6: data <= 32'hEFBF0220;	14'h1FE7: data <= 32'hEFABAE0E;	14'h1FE8: data <= 32'hEF9859FC;	14'h1FE9: data <= 32'hEF867B44;	14'h1FEA: data <= 32'hEF77A2EA;	14'h1FEB: data <= 32'hEF68CA90;	14'h1FEC: data <= 32'hEF59F236;	14'h1FED: data <= 32'hEF4B19DD;	14'h1FEE: data <= 32'hEF3C4183;	14'h1FEF: data <= 32'hEF2D6929;	14'h1FF0: data <= 32'hEF1E90CF;	14'h1FF1: data <= 32'hEF0FB875;	14'h1FF2: data <= 32'hEF00E01B;	14'h1FF3: data <= 32'hEEF207C1;	14'h1FF4: data <= 32'hEEE32F67;	14'h1FF5: data <= 32'hEED4570D;	14'h1FF6: data <= 32'hEEC57EB3;	14'h1FF7: data <= 32'hEEB6A659;	14'h1FF8: data <= 32'hEEA7CDFF;	14'h1FF9: data <= 32'hEE98F5A5;	14'h1FFA: data <= 32'hEE8A1D4C;	14'h1FFB: data <= 32'hEE7B44F2;	14'h1FFC: data <= 32'hEE6C6C98;	14'h1FFD: data <= 32'hEE5D943E;	14'h1FFE: data <= 32'hEE4EBBE4;	14'h1FFF: data <= 32'hEE3FE38A;	14'h2000: data <= 32'hEE310B30;	14'h2001: data <= 32'hEE2232D6;	14'h2002: data <= 32'hEE135A7C;	14'h2003: data <= 32'hEE048222;	14'h2004: data <= 32'hEDF5A9C8;	14'h2005: data <= 32'hEDE6D16E;	14'h2006: data <= 32'hEDD7F914;	14'h2007: data <= 32'hEDC920BB;	14'h2008: data <= 32'hEDBA4861;	14'h2009: data <= 32'hEDAB7007;	14'h200A: data <= 32'hED9C97AD;	14'h200B: data <= 32'hED8DBF53;	14'h200C: data <= 32'hED7EE6F9;	14'h200D: data <= 32'hED711D2E;	14'h200E: data <= 32'hED681DEB;	14'h200F: data <= 32'hED5F1EA8;	14'h2010: data <= 32'hED561F65;	14'h2011: data <= 32'hED4D2022;	14'h2012: data <= 32'hED4420DF;	14'h2013: data <= 32'hED3B219C;	14'h2014: data <= 32'hED322259;	14'h2015: data <= 32'hED292316;	14'h2016: data <= 32'hED2023D3;	14'h2017: data <= 32'hED172490;	14'h2018: data <= 32'hED0E254D;	14'h2019: data <= 32'hED05260A;	14'h201A: data <= 32'hECFC26C7;	14'h201B: data <= 32'hECF32785;	14'h201C: data <= 32'hECEA2842;	14'h201D: data <= 32'hECE128FF;	14'h201E: data <= 32'hECD829BC;	14'h201F: data <= 32'hECCF2A79;	14'h2020: data <= 32'hECC62B36;	14'h2021: data <= 32'hECBD2BF3;	14'h2022: data <= 32'hECB42CB0;	14'h2023: data <= 32'hECAB2D6D;	14'h2024: data <= 32'hECA22E2A;	14'h2025: data <= 32'hEC992EE7;	14'h2026: data <= 32'hEC902FA4;	14'h2027: data <= 32'hEC873061;	14'h2028: data <= 32'hEC7E311E;	14'h2029: data <= 32'hEC7531DB;	14'h202A: data <= 32'hEC6C3298;	14'h202B: data <= 32'hEC633355;	14'h202C: data <= 32'hEC5A3412;	14'h202D: data <= 32'hEC5134CF;	14'h202E: data <= 32'hEC48358C;	14'h202F: data <= 32'hEC3F3649;	14'h2030: data <= 32'hEC363706;	14'h2031: data <= 32'hEC2D87FD;	14'h2032: data <= 32'hEC2D343C;	14'h2033: data <= 32'hEC2CE07C;	14'h2034: data <= 32'hEC2C8CBC;	14'h2035: data <= 32'hEC2C38FC;	14'h2036: data <= 32'hEC2BE53B;	14'h2037: data <= 32'hEC2B917B;	14'h2038: data <= 32'hEC2B3DBB;	14'h2039: data <= 32'hEC2AE9FB;	14'h203A: data <= 32'hEC2A963A;	14'h203B: data <= 32'hEC2A427A;	14'h203C: data <= 32'hEC29EEBA;	14'h203D: data <= 32'hEC299AF9;	14'h203E: data <= 32'hEC294739;	14'h203F: data <= 32'hEC28F379;	14'h2040: data <= 32'hEC289FB9;	14'h2041: data <= 32'hEC284BF8;	14'h2042: data <= 32'hEC27F838;	14'h2043: data <= 32'hEC27A478;	14'h2044: data <= 32'hEC2750B8;	14'h2045: data <= 32'hEC26FCF7;	14'h2046: data <= 32'hEC26A937;	14'h2047: data <= 32'hEC265577;	14'h2048: data <= 32'hEC2601B7;	14'h2049: data <= 32'hEC25ADF6;	14'h204A: data <= 32'hEC255A36;	14'h204B: data <= 32'hEC250676;	14'h204C: data <= 32'hEC24B2B6;	14'h204D: data <= 32'hEC245EF5;	14'h204E: data <= 32'hEC240B35;	14'h204F: data <= 32'hEC23B775;	14'h2050: data <= 32'hEC2363B5;	14'h2051: data <= 32'hEC230FF4;	14'h2052: data <= 32'hEC22BC34;	14'h2053: data <= 32'hEC226874;	14'h2054: data <= 32'hEC2214B4;	14'h2055: data <= 32'hEC21C0F3;	14'h2056: data <= 32'hEC1F6606;	14'h2057: data <= 32'hEC1CCBF4;	14'h2058: data <= 32'hEC1A31E3;	14'h2059: data <= 32'hEC1797D1;	14'h205A: data <= 32'hEC14FDBF;	14'h205B: data <= 32'hEC1263AD;	14'h205C: data <= 32'hEC0FC99B;	14'h205D: data <= 32'hEC0D2F8A;	14'h205E: data <= 32'hEC0A9578;	14'h205F: data <= 32'hEC07FB66;	14'h2060: data <= 32'hEC056154;	14'h2061: data <= 32'hEC02C742;	14'h2062: data <= 32'hEC002D31;	14'h2063: data <= 32'hEBFD931F;	14'h2064: data <= 32'hEBFAF90D;	14'h2065: data <= 32'hEBF85EFB;	14'h2066: data <= 32'hEBF5C4EA;	14'h2067: data <= 32'hEBF32AD8;	14'h2068: data <= 32'hEBF090C6;	14'h2069: data <= 32'hEBEDF6B4;	14'h206A: data <= 32'hEBEB5CA2;	14'h206B: data <= 32'hEBE8C291;	14'h206C: data <= 32'hEBE6287F;	14'h206D: data <= 32'hEBE38E6D;	14'h206E: data <= 32'hEBE0F45B;	14'h206F: data <= 32'hEBDE5A49;	14'h2070: data <= 32'hEBDBC038;	14'h2071: data <= 32'hEBD92626;	14'h2072: data <= 32'hEBD68C14;	14'h2073: data <= 32'hEBD3F202;	14'h2074: data <= 32'hEBD157F0;	14'h2075: data <= 32'hEBCEBDDF;	14'h2076: data <= 32'hEBCC23CD;	14'h2077: data <= 32'hEBC989BB;	14'h2078: data <= 32'hEBC6EFA9;	14'h2079: data <= 32'hEBC45598;	14'h207A: data <= 32'hEBBB1864;	14'h207B: data <= 32'hEBAF9BAE;	14'h207C: data <= 32'hEBA41EF8;	14'h207D: data <= 32'hEB98A242;	14'h207E: data <= 32'hEB8D258C;	14'h207F: data <= 32'hEB81A8D6;	14'h2080: data <= 32'hEB762C1F;	14'h2081: data <= 32'hEB6AAF69;	14'h2082: data <= 32'hEB5F32B3;	14'h2083: data <= 32'hEB53B5FD;	14'h2084: data <= 32'hEB483947;	14'h2085: data <= 32'hEB3CBC90;	14'h2086: data <= 32'hEB313FDA;	14'h2087: data <= 32'hEB25C324;	14'h2088: data <= 32'hEB1A466E;	14'h2089: data <= 32'hEB0EC9B8;	14'h208A: data <= 32'hEB034D02;	14'h208B: data <= 32'hEAF7D04B;	14'h208C: data <= 32'hEAEC5395;	14'h208D: data <= 32'hEAE0D6DF;	14'h208E: data <= 32'hEAD55A29;	14'h208F: data <= 32'hEAC9DD73;	14'h2090: data <= 32'hEABE60BD;	14'h2091: data <= 32'hEAB2E406;	14'h2092: data <= 32'hEAA76750;	14'h2093: data <= 32'hEA9BEA9A;	14'h2094: data <= 32'hEA906DE4;	14'h2095: data <= 32'hEA84F12E;	14'h2096: data <= 32'hEA797478;	14'h2097: data <= 32'hEA6DF7C1;	14'h2098: data <= 32'hEA627B0B;	14'h2099: data <= 32'hEA56FE55;	14'h209A: data <= 32'hEA4B819F;	14'h209B: data <= 32'hEA4004E9;	14'h209C: data <= 32'hEA348833;	14'h209D: data <= 32'hEA290B7C;	14'h209E: data <= 32'hEA155300;	14'h209F: data <= 32'hE9FC2B63;	14'h20A0: data <= 32'hE9E303C5;	14'h20A1: data <= 32'hE9C9DC28;	14'h20A2: data <= 32'hE9B0B48B;	14'h20A3: data <= 32'hE9978CED;	14'h20A4: data <= 32'hE97E6550;	14'h20A5: data <= 32'hE9653DB2;	14'h20A6: data <= 32'hE94C1615;	14'h20A7: data <= 32'hE932EE78;	14'h20A8: data <= 32'hE919C6DA;	14'h20A9: data <= 32'hE9009F3D;	14'h20AA: data <= 32'hE8E7779F;	14'h20AB: data <= 32'hE8CE5002;	14'h20AC: data <= 32'hE8B52865;	14'h20AD: data <= 32'hE89C00C7;	14'h20AE: data <= 32'hE882D92A;	14'h20AF: data <= 32'hE869B18C;	14'h20B0: data <= 32'hE85089EF;	14'h20B1: data <= 32'hE8376252;	14'h20B2: data <= 32'hE81E3AB4;	14'h20B3: data <= 32'hE8051317;	14'h20B4: data <= 32'hE7EBEB79;	14'h20B5: data <= 32'hE7D2C3DC;	14'h20B6: data <= 32'hE7B99C3E;	14'h20B7: data <= 32'hE7A074A1;	14'h20B8: data <= 32'hE7874D04;	14'h20B9: data <= 32'hE76E2566;	14'h20BA: data <= 32'hE754FDC9;	14'h20BB: data <= 32'hE73BD62B;	14'h20BC: data <= 32'hE722AE8E;	14'h20BD: data <= 32'hE70986F1;	14'h20BE: data <= 32'hE6F05F53;	14'h20BF: data <= 32'hE6D737B6;	14'h20C0: data <= 32'hE6BE1018;	14'h20C1: data <= 32'hE6A4E87B;	14'h20C2: data <= 32'hE686E048;	14'h20C3: data <= 32'hE663117E;	14'h20C4: data <= 32'hE63F42B3;	14'h20C5: data <= 32'hE61B73E9;	14'h20C6: data <= 32'hE5F7A51F;	14'h20C7: data <= 32'hE5D3D655;	14'h20C8: data <= 32'hE5B0078B;	14'h20C9: data <= 32'hE58C38C1;	14'h20CA: data <= 32'hE56869F7;	14'h20CB: data <= 32'hE5449B2D;	14'h20CC: data <= 32'hE520CC63;	14'h20CD: data <= 32'hE4FCFD99;	14'h20CE: data <= 32'hE4D92ECE;	14'h20CF: data <= 32'hE4B56004;	14'h20D0: data <= 32'hE491913A;	14'h20D1: data <= 32'hE46DC270;	14'h20D2: data <= 32'hE449F3A6;	14'h20D3: data <= 32'hE42624DC;	14'h20D4: data <= 32'hE4025612;	14'h20D5: data <= 32'hE3DE8748;	14'h20D6: data <= 32'hE3BAB87E;	14'h20D7: data <= 32'hE396E9B4;	14'h20D8: data <= 32'hE3731AEA;	14'h20D9: data <= 32'hE34F4C1F;	14'h20DA: data <= 32'hE32B7D55;	14'h20DB: data <= 32'hE307AE8B;	14'h20DC: data <= 32'hE2E3DFC1;	14'h20DD: data <= 32'hE2C010F7;	14'h20DE: data <= 32'hE29C422D;	14'h20DF: data <= 32'hE2787363;	14'h20E0: data <= 32'hE254A499;	14'h20E1: data <= 32'hE230D5CF;	14'h20E2: data <= 32'hE20D0705;	14'h20E3: data <= 32'hE1E9383B;	14'h20E4: data <= 32'hE1C56970;	14'h20E5: data <= 32'hE1A19AA6;	14'h20E6: data <= 32'hE179A39D;	14'h20E7: data <= 32'hE1488F6C;	14'h20E8: data <= 32'hE1177B3A;	14'h20E9: data <= 32'hE0E66709;	14'h20EA: data <= 32'hE0B552D7;	14'h20EB: data <= 32'hE0843EA6;	14'h20EC: data <= 32'hE0532A74;	14'h20ED: data <= 32'hE0221643;	14'h20EE: data <= 32'hDFF10212;	14'h20EF: data <= 32'hDFBFEDE0;	14'h20F0: data <= 32'hDF8ED9AF;	14'h20F1: data <= 32'hDF5DC57D;	14'h20F2: data <= 32'hDF2CB14C;	14'h20F3: data <= 32'hDEFB9D1A;	14'h20F4: data <= 32'hDECA88E9;	14'h20F5: data <= 32'hDE9974B8;	14'h20F6: data <= 32'hDE686086;	14'h20F7: data <= 32'hDE374C55;	14'h20F8: data <= 32'hDE063823;	14'h20F9: data <= 32'hDDD523F2;	14'h20FA: data <= 32'hDDA40FC0;	14'h20FB: data <= 32'hDD72FB8F;	14'h20FC: data <= 32'hDD41E75E;	14'h20FD: data <= 32'hDD10D32C;	14'h20FE: data <= 32'hDCDFBEFB;	14'h20FF: data <= 32'hDCAEAAC9;	14'h2100: data <= 32'hDC7D9698;	14'h2101: data <= 32'hDC4C8266;	14'h2102: data <= 32'hDC1B6E35;	14'h2103: data <= 32'hDBEA5A04;	14'h2104: data <= 32'hDBB945D2;	14'h2105: data <= 32'hDB8831A1;	14'h2106: data <= 32'hDB571D6F;	14'h2107: data <= 32'hDB26093E;	14'h2108: data <= 32'hDAF4F50C;	14'h2109: data <= 32'hDAC3E0DB;	14'h210A: data <= 32'hDA90433B;	14'h210B: data <= 32'hDA5024D2;	14'h210C: data <= 32'hDA10066A;	14'h210D: data <= 32'hD9CFE802;	14'h210E: data <= 32'hD98FC99A;	14'h210F: data <= 32'hD94FAB32;	14'h2110: data <= 32'hD90F8CCA;	14'h2111: data <= 32'hD8CF6E62;	14'h2112: data <= 32'hD88F4FFA;	14'h2113: data <= 32'hD84F3192;	14'h2114: data <= 32'hD80F1329;	14'h2115: data <= 32'hD7CEF4C1;	14'h2116: data <= 32'hD78ED659;	14'h2117: data <= 32'hD74EB7F1;	14'h2118: data <= 32'hD70E9989;	14'h2119: data <= 32'hD6CE7B21;	14'h211A: data <= 32'hD68E5CB9;	14'h211B: data <= 32'hD64E3E51;	14'h211C: data <= 32'hD60E1FE8;	14'h211D: data <= 32'hD5CE0180;	14'h211E: data <= 32'hD58DE318;	14'h211F: data <= 32'hD54DC4B0;	14'h2120: data <= 32'hD50DA648;	14'h2121: data <= 32'hD4CD87E0;	14'h2122: data <= 32'hD48D6978;	14'h2123: data <= 32'hD44D4B10;	14'h2124: data <= 32'hD40D2CA8;	14'h2125: data <= 32'hD3CD0E3F;	14'h2126: data <= 32'hD38CEFD7;	14'h2127: data <= 32'hD34CD16F;	14'h2128: data <= 32'hD30CB307;	14'h2129: data <= 32'hD2CC949F;	14'h212A: data <= 32'hD28C7637;	14'h212B: data <= 32'hD24C57CF;	14'h212C: data <= 32'hD20C3967;	14'h212D: data <= 32'hD1CC1AFE;	14'h212E: data <= 32'hD18B8944;	14'h212F: data <= 32'hD138B905;	14'h2130: data <= 32'hD0E5E8C6;	14'h2131: data <= 32'hD0931887;	14'h2132: data <= 32'hD0404849;	14'h2133: data <= 32'hCFED780A;	14'h2134: data <= 32'hCF9AA7CB;	14'h2135: data <= 32'hCF47D78C;	14'h2136: data <= 32'hCEF5074D;	14'h2137: data <= 32'hCEA2370E;	14'h2138: data <= 32'hCE4F66CF;	14'h2139: data <= 32'hCDFC9690;	14'h213A: data <= 32'hCDA9C652;	14'h213B: data <= 32'hCD56F613;	14'h213C: data <= 32'hCD0425D4;	14'h213D: data <= 32'hCCB15595;	14'h213E: data <= 32'hCC5E8556;	14'h213F: data <= 32'hCC0BB517;	14'h2140: data <= 32'hCBB8E4D8;	14'h2141: data <= 32'hCB661499;	14'h2142: data <= 32'hCB13445B;	14'h2143: data <= 32'hCAC0741C;	14'h2144: data <= 32'hCA6DA3DD;	14'h2145: data <= 32'hCA1AD39E;	14'h2146: data <= 32'hC9C8035F;	14'h2147: data <= 32'hC9753320;	14'h2148: data <= 32'hC92262E1;	14'h2149: data <= 32'hC8CF92A2;	14'h214A: data <= 32'hC87CC264;	14'h214B: data <= 32'hC829F225;	14'h214C: data <= 32'hC7D721E6;	14'h214D: data <= 32'hC78451A7;	14'h214E: data <= 32'hC7318168;	14'h214F: data <= 32'hC6DEB129;	14'h2150: data <= 32'hC68BE0EA;	14'h2151: data <= 32'hC63910AB;	14'h2152: data <= 32'hC5E6406D;	14'h2153: data <= 32'hC5999D4B;	14'h2154: data <= 32'hC54DD2C1;	14'h2155: data <= 32'hC5020836;	14'h2156: data <= 32'hC4B63DAC;	14'h2157: data <= 32'hC46A7322;	14'h2158: data <= 32'hC41EA898;	14'h2159: data <= 32'hC3D2DE0D;	14'h215A: data <= 32'hC3871383;	14'h215B: data <= 32'hC33B48F9;	14'h215C: data <= 32'hC2EF7E6E;	14'h215D: data <= 32'hC2A3B3E4;	14'h215E: data <= 32'hC257E95A;	14'h215F: data <= 32'hC20C1ED0;	14'h2160: data <= 32'hC1C05445;	14'h2161: data <= 32'hC17489BB;	14'h2162: data <= 32'hC128BF31;	14'h2163: data <= 32'hC0DCF4A6;	14'h2164: data <= 32'hC0912A1C;	14'h2165: data <= 32'hC0455F92;	14'h2166: data <= 32'hBFF99508;	14'h2167: data <= 32'hBFADCA7D;	14'h2168: data <= 32'hBF61FFF3;	14'h2169: data <= 32'hBF163569;	14'h216A: data <= 32'hBECA6ADE;	14'h216B: data <= 32'hBE7EA054;	14'h216C: data <= 32'hBE32D5CA;	14'h216D: data <= 32'hBDE70B40;	14'h216E: data <= 32'hBD9B40B5;	14'h216F: data <= 32'hBD4F762B;	14'h2170: data <= 32'hBD03ABA1;	14'h2171: data <= 32'hBCB7E116;	14'h2172: data <= 32'hBC6C168C;	14'h2173: data <= 32'hBC204C02;	14'h2174: data <= 32'hBBD48178;	14'h2175: data <= 32'hBB88B6ED;	14'h2176: data <= 32'hBB3CEC63;	14'h2177: data <= 32'hBB02B032;	14'h2178: data <= 32'hBACEC8EA;	14'h2179: data <= 32'hBA9AE1A3;	14'h217A: data <= 32'hBA66FA5B;	14'h217B: data <= 32'hBA331313;	14'h217C: data <= 32'hB9FF2BCC;	14'h217D: data <= 32'hB9CB4484;	14'h217E: data <= 32'hB9975D3C;	14'h217F: data <= 32'hB96375F5;	14'h2180: data <= 32'hB92F8EAD;	14'h2181: data <= 32'hB8FBA765;	14'h2182: data <= 32'hB8C7C01E;	14'h2183: data <= 32'hB893D8D6;	14'h2184: data <= 32'hB85FF18E;	14'h2185: data <= 32'hB82C0A47;	14'h2186: data <= 32'hB7F822FF;	14'h2187: data <= 32'hB7C43BB7;	14'h2188: data <= 32'hB7905470;	14'h2189: data <= 32'hB75C6D28;	14'h218A: data <= 32'hB72885E0;	14'h218B: data <= 32'hB6F49E99;	14'h218C: data <= 32'hB6C0B751;	14'h218D: data <= 32'hB68CD009;	14'h218E: data <= 32'hB658E8C2;	14'h218F: data <= 32'hB625017A;	14'h2190: data <= 32'hB5F11A32;	14'h2191: data <= 32'hB5BD32EB;	14'h2192: data <= 32'hB5894BA3;	14'h2193: data <= 32'hB555645C;	14'h2194: data <= 32'hB5217D14;	14'h2195: data <= 32'hB4ED95CC;	14'h2196: data <= 32'hB4B9AE85;	14'h2197: data <= 32'hB485C73D;	14'h2198: data <= 32'hB451DFF5;	14'h2199: data <= 32'hB41DF8AE;	14'h219A: data <= 32'hB3EA1166;	14'h219B: data <= 32'hB377CCD6;	14'h219C: data <= 32'hB2DA4253;	14'h219D: data <= 32'hB23CB7D0;	14'h219E: data <= 32'hB19F2D4D;	14'h219F: data <= 32'hB101A2CA;	14'h21A0: data <= 32'hB0641847;	14'h21A1: data <= 32'hAFC68DC4;	14'h21A2: data <= 32'hAF290341;	14'h21A3: data <= 32'hAE8B78BD;	14'h21A4: data <= 32'hADEDEE3A;	14'h21A5: data <= 32'hAD5063B7;	14'h21A6: data <= 32'hACB2D934;	14'h21A7: data <= 32'hAC154EB1;	14'h21A8: data <= 32'hAB77C42E;	14'h21A9: data <= 32'hAADA39AB;	14'h21AA: data <= 32'hAA3CAF28;	14'h21AB: data <= 32'hA99F24A5;	14'h21AC: data <= 32'hA9019A22;	14'h21AD: data <= 32'hA8640F9F;	14'h21AE: data <= 32'hA7C6851C;	14'h21AF: data <= 32'hA728FA98;	14'h21B0: data <= 32'hA68B7015;	14'h21B1: data <= 32'hA5EDE592;	14'h21B2: data <= 32'hA5505B0F;	14'h21B3: data <= 32'hA4B2D08C;	14'h21B4: data <= 32'hA4154609;	14'h21B5: data <= 32'hA377BB86;	14'h21B6: data <= 32'hA2DA3103;	14'h21B7: data <= 32'hA23CA680;	14'h21B8: data <= 32'hA19F1BFD;	14'h21B9: data <= 32'hA101917A;	14'h21BA: data <= 32'hA06406F6;	14'h21BB: data <= 32'h9FC67C73;	14'h21BC: data <= 32'h9F28F1F0;	14'h21BD: data <= 32'h9E8B676D;	14'h21BE: data <= 32'h9DEDDCEA;	14'h21BF: data <= 32'h9DCB3905;	14'h21C0: data <= 32'h9E4160CE;	14'h21C1: data <= 32'h9EB78898;	14'h21C2: data <= 32'h9F2DB061;	14'h21C3: data <= 32'h9FA3D82A;	14'h21C4: data <= 32'hA019FFF4;	14'h21C5: data <= 32'hA09027BD;	14'h21C6: data <= 32'hA1064F87;	14'h21C7: data <= 32'hA17C7750;	14'h21C8: data <= 32'hA1F29F1A;	14'h21C9: data <= 32'hA268C6E3;	14'h21CA: data <= 32'hA2DEEEAD;	14'h21CB: data <= 32'hA3551676;	14'h21CC: data <= 32'hA3CB3E40;	14'h21CD: data <= 32'hA4416609;	14'h21CE: data <= 32'hA4B78DD3;	14'h21CF: data <= 32'hA52DB59C;	14'h21D0: data <= 32'hA5A3DD66;	14'h21D1: data <= 32'hA61A052F;	14'h21D2: data <= 32'hA6902CF9;	14'h21D3: data <= 32'hA70654C2;	14'h21D4: data <= 32'hA77C7C8C;	14'h21D5: data <= 32'hA7F2A455;	14'h21D6: data <= 32'hA868CC1F;	14'h21D7: data <= 32'hA8DEF3E8;	14'h21D8: data <= 32'hA9551BB2;	14'h21D9: data <= 32'hA9CB437B;	14'h21DA: data <= 32'hAA416B45;	14'h21DB: data <= 32'hAAB7930E;	14'h21DC: data <= 32'hAB2DBAD8;	14'h21DD: data <= 32'hABA3E2A1;	14'h21DE: data <= 32'hAC1A0A6B;	14'h21DF: data <= 32'hAC903234;	14'h21E0: data <= 32'hAD0659FE;	14'h21E1: data <= 32'hAD7C81C7;	14'h21E2: data <= 32'hADF2A990;	14'h21E3: data <= 32'hAE7926C4;	14'h21E4: data <= 32'hAF2588DB;	14'h21E5: data <= 32'hAFD1EAF1;	14'h21E6: data <= 32'hB07E4D07;	14'h21E7: data <= 32'hB12AAF1D;	14'h21E8: data <= 32'hB1D71133;	14'h21E9: data <= 32'hB283734A;	14'h21EA: data <= 32'hB32FD560;	14'h21EB: data <= 32'hB3DC3776;	14'h21EC: data <= 32'hB488998C;	14'h21ED: data <= 32'hB534FBA2;	14'h21EE: data <= 32'hB5E15DB9;	14'h21EF: data <= 32'hB68DBFCF;	14'h21F0: data <= 32'hB73A21E5;	14'h21F1: data <= 32'hB7E683FB;	14'h21F2: data <= 32'hB892E611;	14'h21F3: data <= 32'hB93F4828;	14'h21F4: data <= 32'hB9EBAA3E;	14'h21F5: data <= 32'hBA980C54;	14'h21F6: data <= 32'hBB446E6A;	14'h21F7: data <= 32'hBBF0D080;	14'h21F8: data <= 32'hBC9D3297;	14'h21F9: data <= 32'hBD4994AD;	14'h21FA: data <= 32'hBDF5F6C3;	14'h21FB: data <= 32'hBEA258D9;	14'h21FC: data <= 32'hBF4EBAEF;	14'h21FD: data <= 32'hBFFB1D05;	14'h21FE: data <= 32'hC0A77F1C;	14'h21FF: data <= 32'hC153E132;	14'h2200: data <= 32'hC2004348;	14'h2201: data <= 32'hC2ACA55E;	14'h2202: data <= 32'hC3590774;	14'h2203: data <= 32'hC405698B;	14'h2204: data <= 32'hC4B1CBA1;	14'h2205: data <= 32'hC55E2DB7;	14'h2206: data <= 32'hC60A8FCD;	14'h2207: data <= 32'hC6A69754;	14'h2208: data <= 32'hC6EA8FD5;	14'h2209: data <= 32'hC72E8856;	14'h220A: data <= 32'hC77280D7;	14'h220B: data <= 32'hC7B67958;	14'h220C: data <= 32'hC7FA71DA;	14'h220D: data <= 32'hC83E6A5B;	14'h220E: data <= 32'hC88262DC;	14'h220F: data <= 32'hC8C65B5D;	14'h2210: data <= 32'hC90A53DE;	14'h2211: data <= 32'hC94E4C5F;	14'h2212: data <= 32'hC99244E1;	14'h2213: data <= 32'hC9D63D62;	14'h2214: data <= 32'hCA1A35E3;	14'h2215: data <= 32'hCA5E2E64;	14'h2216: data <= 32'hCAA226E5;	14'h2217: data <= 32'hCAE61F66;	14'h2218: data <= 32'hCB2A17E8;	14'h2219: data <= 32'hCB6E1069;	14'h221A: data <= 32'hCBB208EA;	14'h221B: data <= 32'hCBF6016B;	14'h221C: data <= 32'hCC39F9EC;	14'h221D: data <= 32'hCC7DF26D;	14'h221E: data <= 32'hCCC1EAEE;	14'h221F: data <= 32'hCD05E370;	14'h2220: data <= 32'hCD49DBF1;	14'h2221: data <= 32'hCD8DD472;	14'h2222: data <= 32'hCDD1CCF3;	14'h2223: data <= 32'hCE15C574;	14'h2224: data <= 32'hCE59BDF5;	14'h2225: data <= 32'hCE9DB677;	14'h2226: data <= 32'hCEE1AEF8;	14'h2227: data <= 32'hCF25A779;	14'h2228: data <= 32'hCF699FFA;	14'h2229: data <= 32'hCFAD987B;	14'h222A: data <= 32'hCFF190FC;	14'h222B: data <= 32'hD035223E;	14'h222C: data <= 32'hD057A116;	14'h222D: data <= 32'hD07A1FED;	14'h222E: data <= 32'hD09C9EC5;	14'h222F: data <= 32'hD0BF1D9D;	14'h2230: data <= 32'hD0E19C75;	14'h2231: data <= 32'hD1041B4C;	14'h2232: data <= 32'hD1269A24;	14'h2233: data <= 32'hD14918FC;	14'h2234: data <= 32'hD16B97D4;	14'h2235: data <= 32'hD18E16AB;	14'h2236: data <= 32'hD1B09583;	14'h2237: data <= 32'hD1D3145B;	14'h2238: data <= 32'hD1F59333;	14'h2239: data <= 32'hD218120A;	14'h223A: data <= 32'hD23A90E2;	14'h223B: data <= 32'hD25D0FBA;	14'h223C: data <= 32'hD27F8E92;	14'h223D: data <= 32'hD2A20D6A;	14'h223E: data <= 32'hD2C48C41;	14'h223F: data <= 32'hD2E70B19;	14'h2240: data <= 32'hD30989F1;	14'h2241: data <= 32'hD32C08C9;	14'h2242: data <= 32'hD34E87A0;	14'h2243: data <= 32'hD3710678;	14'h2244: data <= 32'hD3938550;	14'h2245: data <= 32'hD3B60428;	14'h2246: data <= 32'hD3D882FF;	14'h2247: data <= 32'hD3FB01D7;	14'h2248: data <= 32'hD41D80AF;	14'h2249: data <= 32'hD43FFF87;	14'h224A: data <= 32'hD4627E5E;	14'h224B: data <= 32'hD484FD36;	14'h224C: data <= 32'hD4A77C0E;	14'h224D: data <= 32'hD4C9FAE6;	14'h224E: data <= 32'hD4EC79BD;	14'h224F: data <= 32'hD50EF895;	14'h2250: data <= 32'hD523C07C;	14'h2251: data <= 32'hD5366FFF;	14'h2252: data <= 32'hD5491F81;	14'h2253: data <= 32'hD55BCF04;	14'h2254: data <= 32'hD56E7E86;	14'h2255: data <= 32'hD5812E09;	14'h2256: data <= 32'hD593DD8B;	14'h2257: data <= 32'hD5A68D0D;	14'h2258: data <= 32'hD5B93C90;	14'h2259: data <= 32'hD5CBEC12;	14'h225A: data <= 32'hD5DE9B95;	14'h225B: data <= 32'hD5F14B17;	14'h225C: data <= 32'hD603FA9A;	14'h225D: data <= 32'hD616AA1C;	14'h225E: data <= 32'hD629599E;	14'h225F: data <= 32'hD63C0921;	14'h2260: data <= 32'hD64EB8A3;	14'h2261: data <= 32'hD6616826;	14'h2262: data <= 32'hD67417A8;	14'h2263: data <= 32'hD686C72B;	14'h2264: data <= 32'hD69976AD;	14'h2265: data <= 32'hD6AC262F;	14'h2266: data <= 32'hD6BED5B2;	14'h2267: data <= 32'hD6D18534;	14'h2268: data <= 32'hD6E434B7;	14'h2269: data <= 32'hD6F6E439;	14'h226A: data <= 32'hD70993BC;	14'h226B: data <= 32'hD71C433E;	14'h226C: data <= 32'hD72EF2C0;	14'h226D: data <= 32'hD741A243;	14'h226E: data <= 32'hD75451C5;	14'h226F: data <= 32'hD7670148;	14'h2270: data <= 32'hD779B0CA;	14'h2271: data <= 32'hD78C604D;	14'h2272: data <= 32'hD79F0FCF;	14'h2273: data <= 32'hD7B1BF51;	14'h2274: data <= 32'hD7B62F8B;	14'h2275: data <= 32'hD7B529A4;	14'h2276: data <= 32'hD7B423BD;	14'h2277: data <= 32'hD7B31DD6;	14'h2278: data <= 32'hD7B217EF;	14'h2279: data <= 32'hD7B11208;	14'h227A: data <= 32'hD7B00C21;	14'h227B: data <= 32'hD7AF063B;	14'h227C: data <= 32'hD7AE0054;	14'h227D: data <= 32'hD7ACFA6D;	14'h227E: data <= 32'hD7ABF486;	14'h227F: data <= 32'hD7AAEE9F;	14'h2280: data <= 32'hD7A9E8B8;	14'h2281: data <= 32'hD7A8E2D1;	14'h2282: data <= 32'hD7A7DCEA;	14'h2283: data <= 32'hD7A6D703;	14'h2284: data <= 32'hD7A5D11C;	14'h2285: data <= 32'hD7A4CB36;	14'h2286: data <= 32'hD7A3C54F;	14'h2287: data <= 32'hD7A2BF68;	14'h2288: data <= 32'hD7A1B981;	14'h2289: data <= 32'hD7A0B39A;	14'h228A: data <= 32'hD79FADB3;	14'h228B: data <= 32'hD79EA7CC;	14'h228C: data <= 32'hD79DA1E5;	14'h228D: data <= 32'hD79C9BFE;	14'h228E: data <= 32'hD79B9617;	14'h228F: data <= 32'hD79A9031;	14'h2290: data <= 32'hD7998A4A;	14'h2291: data <= 32'hD7988463;	14'h2292: data <= 32'hD7977E7C;	14'h2293: data <= 32'hD7967895;	14'h2294: data <= 32'hD79572AE;	14'h2295: data <= 32'hD7946CC7;	14'h2296: data <= 32'hD79366E0;	14'h2297: data <= 32'hD79260F9;	14'h2298: data <= 32'hD796098C;	14'h2299: data <= 32'hD79D1C02;	14'h229A: data <= 32'hD7A42E79;	14'h229B: data <= 32'hD7AB40EF;	14'h229C: data <= 32'hD7B25366;	14'h229D: data <= 32'hD7B965DC;	14'h229E: data <= 32'hD7C07852;	14'h229F: data <= 32'hD7C78AC9;	14'h22A0: data <= 32'hD7CE9D3F;	14'h22A1: data <= 32'hD7D5AFB5;	14'h22A2: data <= 32'hD7DCC22C;	14'h22A3: data <= 32'hD7E3D4A2;	14'h22A4: data <= 32'hD7EAE718;	14'h22A5: data <= 32'hD7F1F98F;	14'h22A6: data <= 32'hD7F90C05;	14'h22A7: data <= 32'hD8001E7B;	14'h22A8: data <= 32'hD80730F2;	14'h22A9: data <= 32'hD80E4368;	14'h22AA: data <= 32'hD81555DE;	14'h22AB: data <= 32'hD81C6855;	14'h22AC: data <= 32'hD8237ACB;	14'h22AD: data <= 32'hD82A8D41;	14'h22AE: data <= 32'hD8319FB8;	14'h22AF: data <= 32'hD838B22E;	14'h22B0: data <= 32'hD83FC4A4;	14'h22B1: data <= 32'hD846D71B;	14'h22B2: data <= 32'hD84DE991;	14'h22B3: data <= 32'hD854FC07;	14'h22B4: data <= 32'hD85C0E7E;	14'h22B5: data <= 32'hD86320F4;	14'h22B6: data <= 32'hD86A336A;	14'h22B7: data <= 32'hD87145E1;	14'h22B8: data <= 32'hD8785857;	14'h22B9: data <= 32'hD87F6ACD;	14'h22BA: data <= 32'hD8867D44;	14'h22BB: data <= 32'hD88D8FBA;	14'h22BC: data <= 32'hD89C3163;	14'h22BD: data <= 32'hD8B4B18E;	14'h22BE: data <= 32'hD8CD31B9;	14'h22BF: data <= 32'hD8E5B1E4;	14'h22C0: data <= 32'hD8FE320F;	14'h22C1: data <= 32'hD916B23B;	14'h22C2: data <= 32'hD92F3266;	14'h22C3: data <= 32'hD947B291;	14'h22C4: data <= 32'hD96032BC;	14'h22C5: data <= 32'hD978B2E7;	14'h22C6: data <= 32'hD9913312;	14'h22C7: data <= 32'hD9A9B33D;	14'h22C8: data <= 32'hD9C23369;	14'h22C9: data <= 32'hD9DAB394;	14'h22CA: data <= 32'hD9F333BF;	14'h22CB: data <= 32'hDA0BB3EA;	14'h22CC: data <= 32'hDA243415;	14'h22CD: data <= 32'hDA3CB440;	14'h22CE: data <= 32'hDA55346C;	14'h22CF: data <= 32'hDA6DB497;	14'h22D0: data <= 32'hDA8634C2;	14'h22D1: data <= 32'hDA9EB4ED;	14'h22D2: data <= 32'hDAB73518;	14'h22D3: data <= 32'hDACFB543;	14'h22D4: data <= 32'hDAE8356E;	14'h22D5: data <= 32'hDB00B59A;	14'h22D6: data <= 32'hDB1935C5;	14'h22D7: data <= 32'hDB31B5F0;	14'h22D8: data <= 32'hDB4A361B;	14'h22D9: data <= 32'hDB62B646;	14'h22DA: data <= 32'hDB7B3671;	14'h22DB: data <= 32'hDB93B69C;	14'h22DC: data <= 32'hDBAC36C8;	14'h22DD: data <= 32'hDBC4B6F3;	14'h22DE: data <= 32'hDBDD371E;	14'h22DF: data <= 32'hDBF5B749;	14'h22E0: data <= 32'hDC0DB263;	14'h22E1: data <= 32'hDC24665F;	14'h22E2: data <= 32'hDC3B1A5A;	14'h22E3: data <= 32'hDC51CE55;	14'h22E4: data <= 32'hDC688251;	14'h22E5: data <= 32'hDC7F364C;	14'h22E6: data <= 32'hDC95EA48;	14'h22E7: data <= 32'hDCAC9E43;	14'h22E8: data <= 32'hDCC3523E;	14'h22E9: data <= 32'hDCDA063A;	14'h22EA: data <= 32'hDCF0BA35;	14'h22EB: data <= 32'hDD076E31;	14'h22EC: data <= 32'hDD1E222C;	14'h22ED: data <= 32'hDD34D628;	14'h22EE: data <= 32'hDD4B8A23;	14'h22EF: data <= 32'hDD623E1E;	14'h22F0: data <= 32'hDD78F21A;	14'h22F1: data <= 32'hDD8FA615;	14'h22F2: data <= 32'hDDA65A11;	14'h22F3: data <= 32'hDDBD0E0C;	14'h22F4: data <= 32'hDDD3C207;	14'h22F5: data <= 32'hDDEA7603;	14'h22F6: data <= 32'hDE0129FE;	14'h22F7: data <= 32'hDE17DDFA;	14'h22F8: data <= 32'hDE2E91F5;	14'h22F9: data <= 32'hDE4545F0;	14'h22FA: data <= 32'hDE5BF9EC;	14'h22FB: data <= 32'hDE72ADE7;	14'h22FC: data <= 32'hDE8961E3;	14'h22FD: data <= 32'hDEA015DE;	14'h22FE: data <= 32'hDEB6C9D9;	14'h22FF: data <= 32'hDECD7DD5;	14'h2300: data <= 32'hDEE431D0;	14'h2301: data <= 32'hDEFAE5CC;	14'h2302: data <= 32'hDF1199C7;	14'h2303: data <= 32'hDF284DC2;	14'h2304: data <= 32'hDF432944;	14'h2305: data <= 32'hDF76994C;	14'h2306: data <= 32'hDFAA0955;	14'h2307: data <= 32'hDFDD795D;	14'h2308: data <= 32'hE010E965;	14'h2309: data <= 32'hE044596D;	14'h230A: data <= 32'hE077C975;	14'h230B: data <= 32'hE0AB397D;	14'h230C: data <= 32'hE0DEA985;	14'h230D: data <= 32'hE112198E;	14'h230E: data <= 32'hE1458996;	14'h230F: data <= 32'hE178F99E;	14'h2310: data <= 32'hE1AC69A6;	14'h2311: data <= 32'hE1DFD9AE;	14'h2312: data <= 32'hE21349B6;	14'h2313: data <= 32'hE246B9BE;	14'h2314: data <= 32'hE27A29C7;	14'h2315: data <= 32'hE2AD99CF;	14'h2316: data <= 32'hE2E109D7;	14'h2317: data <= 32'hE31479DF;	14'h2318: data <= 32'hE347E9E7;	14'h2319: data <= 32'hE37B59EF;	14'h231A: data <= 32'hE3AEC9F7;	14'h231B: data <= 32'hE3E23A00;	14'h231C: data <= 32'hE415AA08;	14'h231D: data <= 32'hE4491A10;	14'h231E: data <= 32'hE47C8A18;	14'h231F: data <= 32'hE4AFFA20;	14'h2320: data <= 32'hE4E36A28;	14'h2321: data <= 32'hE516DA30;	14'h2322: data <= 32'hE54A4A39;	14'h2323: data <= 32'hE57DBA41;	14'h2324: data <= 32'hE5B12A49;	14'h2325: data <= 32'hE5E49A51;	14'h2326: data <= 32'hE6180A59;	14'h2327: data <= 32'hE64B7A61;	14'h2328: data <= 32'h8A63D707;	14'h2329: data <= 32'h8C5F7ACD;	14'h232A: data <= 32'h8E5B1E92;	14'h232B: data <= 32'h9056C258;	14'h232C: data <= 32'h9252661D;	14'h232D: data <= 32'h944E09E2;	14'h232E: data <= 32'h9649ADA8;	14'h232F: data <= 32'h9845516D;	14'h2330: data <= 32'h9A40F532;	14'h2331: data <= 32'h9C3C98F8;	14'h2332: data <= 32'h9E383CBD;	14'h2333: data <= 32'hA033E082;	14'h2334: data <= 32'hA22F8448;	14'h2335: data <= 32'hA42B280D;	14'h2336: data <= 32'hA626CBD2;	14'h2337: data <= 32'hA8226F98;	14'h2338: data <= 32'hAA1E135D;	14'h2339: data <= 32'hAB2DE45D;	14'h233A: data <= 32'hABFCA75B;	14'h233B: data <= 32'hACCB6A59;	14'h233C: data <= 32'hAD9A2D57;	14'h233D: data <= 32'hAE68F055;	14'h233E: data <= 32'hAF37B353;	14'h233F: data <= 32'hB0067651;	14'h2340: data <= 32'hB0D5394F;	14'h2341: data <= 32'hB1A3FC4D;	14'h2342: data <= 32'hB272BF4B;	14'h2343: data <= 32'hB3418249;	14'h2344: data <= 32'hB4104547;	14'h2345: data <= 32'hB4DF0845;	14'h2346: data <= 32'hB5ADCB43;	14'h2347: data <= 32'hB67C8E41;	14'h2348: data <= 32'hB74B513F;	14'h2349: data <= 32'hB7D6723E;	14'h234A: data <= 32'hB82E0BA1;	14'h234B: data <= 32'hB885A504;	14'h234C: data <= 32'hB8DD3E67;	14'h234D: data <= 32'hB934D7CA;	14'h234E: data <= 32'hB98C712C;	14'h234F: data <= 32'hB9E40A8F;	14'h2350: data <= 32'hBA3BA3F2;	14'h2351: data <= 32'hBA933D55;	14'h2352: data <= 32'hBAEAD6B8;	14'h2353: data <= 32'hBB42701A;	14'h2354: data <= 32'hBB9A097D;	14'h2355: data <= 32'hBBF1A2E0;	14'h2356: data <= 32'hBC493C43;	14'h2357: data <= 32'hBCA0D5A5;	14'h2358: data <= 32'hBCF86F08;	14'h2359: data <= 32'hBD49BB61;	14'h235A: data <= 32'hBD8F65CE;	14'h235B: data <= 32'hBDD5103C;	14'h235C: data <= 32'hBE1ABAA9;	14'h235D: data <= 32'hBE606517;	14'h235E: data <= 32'hBEA60F84;	14'h235F: data <= 32'hBEEBB9F2;	14'h2360: data <= 32'hBF31645F;	14'h2361: data <= 32'hBF770ECD;	14'h2362: data <= 32'hBFBCB93A;	14'h2363: data <= 32'hC00263A8;	14'h2364: data <= 32'hC0480E15;	14'h2365: data <= 32'hC08DB882;	14'h2366: data <= 32'hC0D362F0;	14'h2367: data <= 32'hC1190D5D;	14'h2368: data <= 32'hC15EB7CB;	14'h2369: data <= 32'hC1A72E7B;	14'h236A: data <= 32'hC2018D3C;	14'h236B: data <= 32'hC25BEBFD;	14'h236C: data <= 32'hC2B64ABF;	14'h236D: data <= 32'hC310A980;	14'h236E: data <= 32'hC36B0841;	14'h236F: data <= 32'hC3C56702;	14'h2370: data <= 32'hC41FC5C3;	14'h2371: data <= 32'hC47A2484;	14'h2372: data <= 32'hC4D48346;	14'h2373: data <= 32'hC52EE207;	14'h2374: data <= 32'hC58940C8;	14'h2375: data <= 32'hC5E39F89;	14'h2376: data <= 32'hC63DFE4A;	14'h2377: data <= 32'hC6985D0C;	14'h2378: data <= 32'hC6F2BBCD;	14'h2379: data <= 32'hC74D1A8E;	14'h237A: data <= 32'hC7A617AA;	14'h237B: data <= 32'hC7FEF591;	14'h237C: data <= 32'hC857D379;	14'h237D: data <= 32'hC8B0B161;	14'h237E: data <= 32'hC9098F48;	14'h237F: data <= 32'hC9626D30;	14'h2380: data <= 32'hC9BB4B17;	14'h2381: data <= 32'hCA1428FF;	14'h2382: data <= 32'hCA6D06E6;	14'h2383: data <= 32'hCAC5E4CE;	14'h2384: data <= 32'hCB1EC2B5;	14'h2385: data <= 32'hCB77A09D;	14'h2386: data <= 32'hCBD07E85;	14'h2387: data <= 32'hCC295C6C;	14'h2388: data <= 32'hCC823A54;	14'h2389: data <= 32'hCCDB183B;	14'h238A: data <= 32'hCD164E43;	14'h238B: data <= 32'hCD44F858;	14'h238C: data <= 32'hCD73A26D;	14'h238D: data <= 32'hCDA24C82;	14'h238E: data <= 32'hCDD0F697;	14'h238F: data <= 32'hCDFFA0AD;	14'h2390: data <= 32'hCE2E4AC2;	14'h2391: data <= 32'hCE5CF4D7;	14'h2392: data <= 32'hCE8B9EEC;	14'h2393: data <= 32'hCEBA4901;	14'h2394: data <= 32'hCEE8F316;	14'h2395: data <= 32'hCF179D2B;	14'h2396: data <= 32'hCF464741;	14'h2397: data <= 32'hCF74F156;	14'h2398: data <= 32'hCFA39B6B;	14'h2399: data <= 32'hCFD24580;	14'h239A: data <= 32'hCFF05940;	14'h239B: data <= 32'hCFFCEAC3;	14'h239C: data <= 32'hD0097C47;	14'h239D: data <= 32'hD0160DCA;	14'h239E: data <= 32'hD0229F4D;	14'h239F: data <= 32'hD02F30D0;	14'h23A0: data <= 32'hD03BC253;	14'h23A1: data <= 32'hD04853D6;	14'h23A2: data <= 32'hD054E559;	14'h23A3: data <= 32'hD06176DD;	14'h23A4: data <= 32'hD06E0860;	14'h23A5: data <= 32'hD07A99E3;	14'h23A6: data <= 32'hD0872B66;	14'h23A7: data <= 32'hD093BCE9;	14'h23A8: data <= 32'hD0A04E6C;	14'h23A9: data <= 32'hD0ACDFEF;	14'h23AA: data <= 32'hD0BAED32;	14'h23AB: data <= 32'hD0CCFBC8;	14'h23AC: data <= 32'hD0DF0A5E;	14'h23AD: data <= 32'hD0F118F4;	14'h23AE: data <= 32'hD103278A;	14'h23AF: data <= 32'hD115361F;	14'h23B0: data <= 32'hD12744B5;	14'h23B1: data <= 32'hD139534B;	14'h23B2: data <= 32'hD14B61E1;	14'h23B3: data <= 32'hD15D7077;	14'h23B4: data <= 32'hD16F7F0C;	14'h23B5: data <= 32'hD1818DA2;	14'h23B6: data <= 32'hD1939C38;	14'h23B7: data <= 32'hD1A5AACE;	14'h23B8: data <= 32'hD1B7B963;	14'h23B9: data <= 32'hD1C9C7F9;	14'h23BA: data <= 32'hD1DCB3F4;	14'h23BB: data <= 32'hD1FEC24B;	14'h23BC: data <= 32'hD220D0A3;	14'h23BD: data <= 32'hD242DEFB;	14'h23BE: data <= 32'hD264ED53;	14'h23BF: data <= 32'hD286FBAB;	14'h23C0: data <= 32'hD2A90A02;	14'h23C1: data <= 32'hD2CB185A;	14'h23C2: data <= 32'hD2ED26B2;	14'h23C3: data <= 32'hD30F350A;	14'h23C4: data <= 32'hD3314362;	14'h23C5: data <= 32'hD35351B9;	14'h23C6: data <= 32'hD3756011;	14'h23C7: data <= 32'hD3976E69;	14'h23C8: data <= 32'hD3B97CC1;	14'h23C9: data <= 32'hD3DB8B19;	14'h23CA: data <= 32'hD3FD9970;	14'h23CB: data <= 32'hD4225872;	14'h23CC: data <= 32'hD4479CBE;	14'h23CD: data <= 32'hD46CE10A;	14'h23CE: data <= 32'hD4922556;	14'h23CF: data <= 32'hD4B769A2;	14'h23D0: data <= 32'hD4DCADEE;	14'h23D1: data <= 32'hD501F23A;	14'h23D2: data <= 32'hD5273686;	14'h23D3: data <= 32'hD54C7AD2;	14'h23D4: data <= 32'hD571BF1D;	14'h23D5: data <= 32'hD5970369;	14'h23D6: data <= 32'hD5BC47B5;	14'h23D7: data <= 32'hD5E18C01;	14'h23D8: data <= 32'hD606D04D;	14'h23D9: data <= 32'hD62C1499;	14'h23DA: data <= 32'hD65158E5;	14'h23DB: data <= 32'hD674FA75;	14'h23DC: data <= 32'hD6979D23;	14'h23DD: data <= 32'hD6BA3FD1;	14'h23DE: data <= 32'hD6DCE27F;	14'h23DF: data <= 32'hD6FF852D;	14'h23E0: data <= 32'hD72227DB;	14'h23E1: data <= 32'hD744CA88;	14'h23E2: data <= 32'hD7676D36;	14'h23E3: data <= 32'hD78A0FE4;	14'h23E4: data <= 32'hD7ACB292;	14'h23E5: data <= 32'hD7CF5540;	14'h23E6: data <= 32'hD7F1F7EE;	14'h23E7: data <= 32'hD8149A9C;	14'h23E8: data <= 32'hD8373D4A;	14'h23E9: data <= 32'hD859DFF8;	14'h23EA: data <= 32'hD87C82A6;	14'h23EB: data <= 32'hD89E0971;	14'h23EC: data <= 32'hD8BDEFDC;	14'h23ED: data <= 32'hD8DDD648;	14'h23EE: data <= 32'hD8FDBCB4;	14'h23EF: data <= 32'hD91DA31F;	14'h23F0: data <= 32'hD93D898B;	14'h23F1: data <= 32'hD95D6FF7;	14'h23F2: data <= 32'hD97D5663;	14'h23F3: data <= 32'hD99D3CCE;	14'h23F4: data <= 32'hD9BD233A;	14'h23F5: data <= 32'hD9DD09A6;	14'h23F6: data <= 32'hD9FCF012;	14'h23F7: data <= 32'hDA1CD67D;	14'h23F8: data <= 32'hDA3CBCE9;	14'h23F9: data <= 32'hDA5CA355;	14'h23FA: data <= 32'hDA7C89C0;	14'h23FB: data <= 32'hDA9A13C7;	14'h23FC: data <= 32'hDAAD7F8C;	14'h23FD: data <= 32'hDAC0EB51;	14'h23FE: data <= 32'hDAD45716;	14'h23FF: data <= 32'hDAE7C2DB;	14'h2400: data <= 32'hDAFB2EA0;	14'h2401: data <= 32'hDB0E9A65;	14'h2402: data <= 32'hDB22062A;	14'h2403: data <= 32'hDB3571EF;	14'h2404: data <= 32'hDB48DDB4;	14'h2405: data <= 32'hDB5C4979;	14'h2406: data <= 32'hDB6FB53E;	14'h2407: data <= 32'hDB832103;	14'h2408: data <= 32'hDB968CC7;	14'h2409: data <= 32'hDBA9F88C;	14'h240A: data <= 32'hDBBD6451;	14'h240B: data <= 32'hDBD0D016;	14'h240C: data <= 32'hDBDB34DC;	14'h240D: data <= 32'hDBE55970;	14'h240E: data <= 32'hDBEF7E04;	14'h240F: data <= 32'hDBF9A298;	14'h2410: data <= 32'hDC03C72C;	14'h2411: data <= 32'hDC0DEBC0;	14'h2412: data <= 32'hDC181054;	14'h2413: data <= 32'hDC2234E8;	14'h2414: data <= 32'hDC2C597C;	14'h2415: data <= 32'hDC367E11;	14'h2416: data <= 32'hDC40A2A5;	14'h2417: data <= 32'hDC4AC739;	14'h2418: data <= 32'hDC54EBCD;	14'h2419: data <= 32'hDC5F1061;	14'h241A: data <= 32'hDC6934F5;	14'h241B: data <= 32'hDC735989;	14'h241C: data <= 32'hDC7BAEDA;	14'h241D: data <= 32'hDC836F43;	14'h241E: data <= 32'hDC8B2FAC;	14'h241F: data <= 32'hDC92F015;	14'h2420: data <= 32'hDC9AB07E;	14'h2421: data <= 32'hDCA270E7;	14'h2422: data <= 32'hDCAA3150;	14'h2423: data <= 32'hDCB1F1B9;	14'h2424: data <= 32'hDCB9B222;	14'h2425: data <= 32'hDCC1728B;	14'h2426: data <= 32'hDCC932F5;	14'h2427: data <= 32'hDCD0F35E;	14'h2428: data <= 32'hDCD8B3C7;	14'h2429: data <= 32'hDCE07430;	14'h242A: data <= 32'hDCE83499;	14'h242B: data <= 32'hDCEFF502;	14'h242C: data <= 32'hDCF37158;	14'h242D: data <= 32'hDCF34D6C;	14'h242E: data <= 32'hDCF3297F;	14'h242F: data <= 32'hDCF30593;	14'h2430: data <= 32'hDCF2E1A7;	14'h2431: data <= 32'hDCF2BDBA;	14'h2432: data <= 32'hDCF299CE;	14'h2433: data <= 32'hDCF275E1;	14'h2434: data <= 32'hDCF251F5;	14'h2435: data <= 32'hDCF22E08;	14'h2436: data <= 32'hDCF20A1C;	14'h2437: data <= 32'hDCF1E62F;	14'h2438: data <= 32'hDCF1C243;	14'h2439: data <= 32'hDCF19E56;	14'h243A: data <= 32'hDCF17A6A;	14'h243B: data <= 32'hDCF1567D;	14'h243C: data <= 32'hDCEEF71C;	14'h243D: data <= 32'hDCE7F132;	14'h243E: data <= 32'hDCE0EB47;	14'h243F: data <= 32'hDCD9E55D;	14'h2440: data <= 32'hDCD2DF72;	14'h2441: data <= 32'hDCCBD988;	14'h2442: data <= 32'hDCC4D39E;	14'h2443: data <= 32'hDCBDCDB3;	14'h2444: data <= 32'hDCB6C7C9;	14'h2445: data <= 32'hDCAFC1DF;	14'h2446: data <= 32'hDCA8BBF4;	14'h2447: data <= 32'hDCA1B60A;	14'h2448: data <= 32'hDC9AB01F;	14'h2449: data <= 32'hDC93AA35;	14'h244A: data <= 32'hDC8CA44B;	14'h244B: data <= 32'hDC859E60;	14'h244C: data <= 32'hDC7EDF13;	14'h244D: data <= 32'hDC7A6652;	14'h244E: data <= 32'hDC75ED91;	14'h244F: data <= 32'hDC7174D0;	14'h2450: data <= 32'hDC6CFC10;	14'h2451: data <= 32'hDC68834F;	14'h2452: data <= 32'hDC640A8E;	14'h2453: data <= 32'hDC5F91CD;	14'h2454: data <= 32'hDC5B190C;	14'h2455: data <= 32'hDC56A04C;	14'h2456: data <= 32'hDC52278B;	14'h2457: data <= 32'hDC4DAECA;	14'h2458: data <= 32'hDC493609;	14'h2459: data <= 32'hDC44BD49;	14'h245A: data <= 32'hDC404488;	14'h245B: data <= 32'hDC3BCBC7;	14'h245C: data <= 32'hDC375306;	14'h245D: data <= 32'hDC383180;	14'h245E: data <= 32'hDC39B5B4;	14'h245F: data <= 32'hDC3B39E8;	14'h2460: data <= 32'hDC3CBE1B;	14'h2461: data <= 32'hDC3E424F;	14'h2462: data <= 32'hDC3FC683;	14'h2463: data <= 32'hDC414AB6;	14'h2464: data <= 32'hDC42CEEA;	14'h2465: data <= 32'hDC44531E;	14'h2466: data <= 32'hDC45D751;	14'h2467: data <= 32'hDC475B85;	14'h2468: data <= 32'hDC48DFB9;	14'h2469: data <= 32'hDC4A63EC;	14'h246A: data <= 32'hDC4BE820;	14'h246B: data <= 32'hDC4D6C54;	14'h246C: data <= 32'hDC4EF087;	14'h246D: data <= 32'hDC56395F;	14'h246E: data <= 32'hDC604701;	14'h246F: data <= 32'hDC6A54A3;	14'h2470: data <= 32'hDC746244;	14'h2471: data <= 32'hDC7E6FE6;	14'h2472: data <= 32'hDC887D88;	14'h2473: data <= 32'hDC928B2A;	14'h2474: data <= 32'hDC9C98CB;	14'h2475: data <= 32'hDCA6A66D;	14'h2476: data <= 32'hDCB0B40F;	14'h2477: data <= 32'hDCBAC1B1;	14'h2478: data <= 32'hDCC4CF52;	14'h2479: data <= 32'hDCCEDCF4;	14'h247A: data <= 32'hDCD8EA96;	14'h247B: data <= 32'hDCE2F838;	14'h247C: data <= 32'hDCED05D9;	14'h247D: data <= 32'hDCF6B069;	14'h247E: data <= 32'hDCFFE669;	14'h247F: data <= 32'hDD091C6A;	14'h2480: data <= 32'hDD12526A;	14'h2481: data <= 32'hDD1B886B;	14'h2482: data <= 32'hDD24BE6B;	14'h2483: data <= 32'hDD2DF46C;	14'h2484: data <= 32'hDD372A6D;	14'h2485: data <= 32'hDD40606D;	14'h2486: data <= 32'hDD49966E;	14'h2487: data <= 32'hDD52CC6E;	14'h2488: data <= 32'hDD5C026F;	14'h2489: data <= 32'hDD653870;	14'h248A: data <= 32'hDD6E6E70;	14'h248B: data <= 32'hDD77A471;	14'h248C: data <= 32'hDD80DA71;	14'h248D: data <= 32'hDD87F277;	14'h248E: data <= 32'hDD887453;	14'h248F: data <= 32'hDD88F62F;	14'h2490: data <= 32'hDD89780A;	14'h2491: data <= 32'hDD89F9E6;	14'h2492: data <= 32'hDD8A7BC2;	14'h2493: data <= 32'hDD8AFD9E;	14'h2494: data <= 32'hDD8B7F7A;	14'h2495: data <= 32'hDD8C0156;	14'h2496: data <= 32'hDD8C8332;	14'h2497: data <= 32'hDD8D050E;	14'h2498: data <= 32'hDD8D86EA;	14'h2499: data <= 32'hDD8E08C5;	14'h249A: data <= 32'hDD8E8AA1;	14'h249B: data <= 32'hDD8F0C7D;	14'h249C: data <= 32'hDD8F8E59;	14'h249D: data <= 32'hDD902304;	14'h249E: data <= 32'hDD935CC0;	14'h249F: data <= 32'hDD96967C;	14'h24A0: data <= 32'hDD99D038;	14'h24A1: data <= 32'hDD9D09F4;	14'h24A2: data <= 32'hDDA043B0;	14'h24A3: data <= 32'hDDA37D6C;	14'h24A4: data <= 32'hDDA6B728;	14'h24A5: data <= 32'hDDA9F0E4;	14'h24A6: data <= 32'hDDAD2AA1;	14'h24A7: data <= 32'hDDB0645D;	14'h24A8: data <= 32'hDDB39E19;	14'h24A9: data <= 32'hDDB6D7D5;	14'h24AA: data <= 32'hDDBA1191;	14'h24AB: data <= 32'hDDBD4B4D;	14'h24AC: data <= 32'hDDC08509;	14'h24AD: data <= 32'hDDC3BEC5;	14'h24AE: data <= 32'hDDC86C0E;	14'h24AF: data <= 32'hDDCD7009;	14'h24B0: data <= 32'hDDD27404;	14'h24B1: data <= 32'hDDD777FE;	14'h24B2: data <= 32'hDDDC7BF9;	14'h24B3: data <= 32'hDDE17FF4;	14'h24B4: data <= 32'hDDE683EF;	14'h24B5: data <= 32'hDDEB87EA;	14'h24B6: data <= 32'hDDF08BE5;	14'h24B7: data <= 32'hDDF58FDF;	14'h24B8: data <= 32'hDDFA93DA;	14'h24B9: data <= 32'hDDFF97D5;	14'h24BA: data <= 32'hDE049BD0;	14'h24BB: data <= 32'hDE099FCB;	14'h24BC: data <= 32'hDE0EA3C5;	14'h24BD: data <= 32'hDE13A7C0;	14'h24BE: data <= 32'hDE180CC1;	14'h24BF: data <= 32'hDE1C055E;	14'h24C0: data <= 32'hDE1FFDFB;	14'h24C1: data <= 32'hDE23F698;	14'h24C2: data <= 32'hDE27EF35;	14'h24C3: data <= 32'hDE2BE7D2;	14'h24C4: data <= 32'hDE2FE06F;	14'h24C5: data <= 32'hDE33D90C;	14'h24C6: data <= 32'hDE37D1A9;	14'h24C7: data <= 32'hDE3BCA46;	14'h24C8: data <= 32'hDE3FC2E3;	14'h24C9: data <= 32'hDE43BB80;	14'h24CA: data <= 32'hDE47B41D;	14'h24CB: data <= 32'hDE4BACBA;	14'h24CC: data <= 32'hDE4FA557;	14'h24CD: data <= 32'hDE539DF4;	14'h24CE: data <= 32'hDE5A6E7F;	14'h24CF: data <= 32'hDE65EAEE;	14'h24D0: data <= 32'hDE71675D;	14'h24D1: data <= 32'hDE7CE3CD;	14'h24D2: data <= 32'hDE88603C;	14'h24D3: data <= 32'hDE93DCAB;	14'h24D4: data <= 32'hDE9F591A;	14'h24D5: data <= 32'hDEAAD589;	14'h24D6: data <= 32'hDEB651F8;	14'h24D7: data <= 32'hDEC1CE67;	14'h24D8: data <= 32'hDECD4AD6;	14'h24D9: data <= 32'hDED8C746;	14'h24DA: data <= 32'hDEE443B5;	14'h24DB: data <= 32'hDEEFC024;	14'h24DC: data <= 32'hDEFB3C93;	14'h24DD: data <= 32'hDF06B902;	14'h24DE: data <= 32'hDF124465;	14'h24DF: data <= 32'hDF1E1D0C;	14'h24E0: data <= 32'hDF29F5B2;	14'h24E1: data <= 32'hDF35CE59;	14'h24E2: data <= 32'hDF41A6FF;	14'h24E3: data <= 32'hDF4D7FA6;	14'h24E4: data <= 32'hDF59584C;	14'h24E5: data <= 32'hDF6530F2;	14'h24E6: data <= 32'hDF710999;	14'h24E7: data <= 32'hDF7CE23F;	14'h24E8: data <= 32'hDF88BAE6;	14'h24E9: data <= 32'hDF94938C;	14'h24EA: data <= 32'hDFA06C32;	14'h24EB: data <= 32'hDFAC44D9;	14'h24EC: data <= 32'hDFB81D7F;	14'h24ED: data <= 32'hDFC3F626;	14'h24EE: data <= 32'hDFCFCECC;	14'h24EF: data <= 32'hDFD60925;	14'h24F0: data <= 32'hDFDBF14D;	14'h24F1: data <= 32'hDFE1D975;	14'h24F2: data <= 32'hDFE7C19D;	14'h24F3: data <= 32'hDFEDA9C5;	14'h24F4: data <= 32'hDFF391EE;	14'h24F5: data <= 32'hDFF97A16;	14'h24F6: data <= 32'hDFFF623E;	14'h24F7: data <= 32'hE0054A66;	14'h24F8: data <= 32'hE00B328E;	14'h24F9: data <= 32'hE0111AB7;	14'h24FA: data <= 32'hE01702DF;	14'h24FB: data <= 32'hE01CEB07;	14'h24FC: data <= 32'hE022D32F;	14'h24FD: data <= 32'hE028BB57;	14'h24FE: data <= 32'hE02EA380;	14'h24FF: data <= 32'hE037355D;	14'h2500: data <= 32'hE040C3B7;	14'h2501: data <= 32'hE04A5211;	14'h2502: data <= 32'hE053E06B;	14'h2503: data <= 32'hE05D6EC5;	14'h2504: data <= 32'hE066FD1F;	14'h2505: data <= 32'hE0708B79;	14'h2506: data <= 32'hE07A19D3;	14'h2507: data <= 32'hE083A82C;	14'h2508: data <= 32'hE08D3686;	14'h2509: data <= 32'hE096C4E0;	14'h250A: data <= 32'hE0A0533A;	14'h250B: data <= 32'hE0A9E194;	14'h250C: data <= 32'hE0B36FEE;	14'h250D: data <= 32'hE0BCFE48;	14'h250E: data <= 32'hE0C68CA2;	14'h250F: data <= 32'hE0D0B6FE;	14'h2510: data <= 32'hE0DB7526;	14'h2511: data <= 32'hE0E6334E;	14'h2512: data <= 32'hE0F0F177;	14'h2513: data <= 32'hE0FBAF9F;	14'h2514: data <= 32'hE1066DC7;	14'h2515: data <= 32'hE1112BF0;	14'h2516: data <= 32'hE11BEA18;	14'h2517: data <= 32'hE126A840;	14'h2518: data <= 32'hE1316669;	14'h2519: data <= 32'hE13C2491;	14'h251A: data <= 32'hE146E2B9;	14'h251B: data <= 32'hE151A0E2;	14'h251C: data <= 32'hE15C5F0A;	14'h251D: data <= 32'hE1671D32;	14'h251E: data <= 32'hE171DB5A;	14'h251F: data <= 32'hE17C41D2;	14'h2520: data <= 32'hE185D906;	14'h2521: data <= 32'hE18F703A;	14'h2522: data <= 32'hE199076E;	14'h2523: data <= 32'hE1A29EA2;	14'h2524: data <= 32'hE1AC35D6;	14'h2525: data <= 32'hE1B5CD0A;	14'h2526: data <= 32'hE1BF643E;	14'h2527: data <= 32'hE1C8FB72;	14'h2528: data <= 32'hE1D292A6;	14'h2529: data <= 32'hE1DC29DA;	14'h252A: data <= 32'hE1E5C10E;	14'h252B: data <= 32'hE1EF5842;	14'h252C: data <= 32'hE1F8EF76;	14'h252D: data <= 32'hE20286AA;	14'h252E: data <= 32'hE20C1DDE;	14'h252F: data <= 32'hE215ACF5;	14'h2530: data <= 32'hE21EE020;	14'h2531: data <= 32'hE228134A;	14'h2532: data <= 32'hE2314675;	14'h2533: data <= 32'hE23A799F;	14'h2534: data <= 32'hE243ACCA;	14'h2535: data <= 32'hE24CDFF4;	14'h2536: data <= 32'hE256131F;	14'h2537: data <= 32'hE25F4649;	14'h2538: data <= 32'hE2687974;	14'h2539: data <= 32'hE271AC9E;	14'h253A: data <= 32'hE27ADFC9;	14'h253B: data <= 32'hE28412F3;	14'h253C: data <= 32'hE28D461E;	14'h253D: data <= 32'hE2967948;	14'h253E: data <= 32'hE29FAC73;	14'h253F: data <= 32'hE2A8DF9D;	14'h2540: data <= 32'hE2B2F094;	14'h2541: data <= 32'hE2BD2432;	14'h2542: data <= 32'hE2C757D1;	14'h2543: data <= 32'hE2D18B6F;	14'h2544: data <= 32'hE2DBBF0D;	14'h2545: data <= 32'hE2E5F2AC;	14'h2546: data <= 32'hE2F0264A;	14'h2547: data <= 32'hE2FA59E8;	14'h2548: data <= 32'hE3048D87;	14'h2549: data <= 32'hE30EC125;	14'h254A: data <= 32'hE318F4C3;	14'h254B: data <= 32'hE3232862;	14'h254C: data <= 32'hE32D5C00;	14'h254D: data <= 32'hE3378F9E;	14'h254E: data <= 32'hE341C33D;	14'h254F: data <= 32'hE34BF6DB;	14'h2550: data <= 32'hE35657BD;	14'h2551: data <= 32'hE360D125;	14'h2552: data <= 32'hE36B4A8C;	14'h2553: data <= 32'hE375C3F3;	14'h2554: data <= 32'hE3803D5B;	14'h2555: data <= 32'hE38AB6C2;	14'h2556: data <= 32'hE3953029;	14'h2557: data <= 32'hE39FA990;	14'h2558: data <= 32'hE3AA22F8;	14'h2559: data <= 32'hE3B49C5F;	14'h255A: data <= 32'hE3BF15C6;	14'h255B: data <= 32'hE3C98F2E;	14'h255C: data <= 32'hE3D40895;	14'h255D: data <= 32'hE3DE81FC;	14'h255E: data <= 32'hE3E8FB64;	14'h255F: data <= 32'hE3F374CB;	14'h2560: data <= 32'hE3FB9A4E;	14'h2561: data <= 32'hE400B1B5;	14'h2562: data <= 32'hE405C91C;	14'h2563: data <= 32'hE40AE083;	14'h2564: data <= 32'hE40FF7EA;	14'h2565: data <= 32'hE4150F51;	14'h2566: data <= 32'hE41A26B8;	14'h2567: data <= 32'hE41F3E20;	14'h2568: data <= 32'hE4245587;	14'h2569: data <= 32'hE4296CEE;	14'h256A: data <= 32'hE42E8455;	14'h256B: data <= 32'hE4339BBC;	14'h256C: data <= 32'hE438B323;	14'h256D: data <= 32'hE43DCA8A;	14'h256E: data <= 32'hE442E1F1;	14'h256F: data <= 32'hE447F958;	14'h2570: data <= 32'hE44B7A90;	14'h2571: data <= 32'hE4493B59;	14'h2572: data <= 32'hE446FC23;	14'h2573: data <= 32'hE444BCEC;	14'h2574: data <= 32'hE4427DB6;	14'h2575: data <= 32'hE4403E7F;	14'h2576: data <= 32'hE43DFF49;	14'h2577: data <= 32'hE43BC013;	14'h2578: data <= 32'hE43980DC;	14'h2579: data <= 32'hE43741A6;	14'h257A: data <= 32'hE435026F;	14'h257B: data <= 32'hE432C339;	14'h257C: data <= 32'hE4308402;	14'h257D: data <= 32'hE42E44CC;	14'h257E: data <= 32'hE42C0595;	14'h257F: data <= 32'hE429C65F;	14'h2580: data <= 32'hE4278728;	14'h2581: data <= 32'hE422FA09;	14'h2582: data <= 32'hE41E6CEA;	14'h2583: data <= 32'hE419DFCB;	14'h2584: data <= 32'hE41552AC;	14'h2585: data <= 32'hE410C58D;	14'h2586: data <= 32'hE40C386E;	14'h2587: data <= 32'hE407AB4F;	14'h2588: data <= 32'hE4031E30;	14'h2589: data <= 32'hE3FE9111;	14'h258A: data <= 32'hE3FA03F2;	14'h258B: data <= 32'hE3F576D3;	14'h258C: data <= 32'hE3F0E9B4;	14'h258D: data <= 32'hE3EC5C95;	14'h258E: data <= 32'hE3E7CF76;	14'h258F: data <= 32'hE3E34257;	14'h2590: data <= 32'hE3DEB538;	14'h2591: data <= 32'hE3DD04A3;	14'h2592: data <= 32'hE3DC1E24;	14'h2593: data <= 32'hE3DB37A5;	14'h2594: data <= 32'hE3DA5125;	14'h2595: data <= 32'hE3D96AA6;	14'h2596: data <= 32'hE3D88426;	14'h2597: data <= 32'hE3D79DA7;	14'h2598: data <= 32'hE3D6B728;	14'h2599: data <= 32'hE3D5D0A8;	14'h259A: data <= 32'hE3D4EA29;	14'h259B: data <= 32'hE3D403A9;	14'h259C: data <= 32'hE3D31D2A;	14'h259D: data <= 32'hE3D236AA;	14'h259E: data <= 32'hE3D1502B;	14'h259F: data <= 32'hE3D069AC;	14'h25A0: data <= 32'hE3CF832C;	14'h25A1: data <= 32'hE3D01719;	14'h25A2: data <= 32'hE3D1CB57;	14'h25A3: data <= 32'hE3D37F95;	14'h25A4: data <= 32'hE3D533D4;	14'h25A5: data <= 32'hE3D6E812;	14'h25A6: data <= 32'hE3D89C51;	14'h25A7: data <= 32'hE3DA508F;	14'h25A8: data <= 32'hE3DC04CD;	14'h25A9: data <= 32'hE3DDB90C;	14'h25AA: data <= 32'hE3DF6D4A;	14'h25AB: data <= 32'hE3E12188;	14'h25AC: data <= 32'hE3E2D5C7;	14'h25AD: data <= 32'hE3E48A05;	14'h25AE: data <= 32'hE3E63E44;	14'h25AF: data <= 32'hE3E7F282;	14'h25B0: data <= 32'hE3E9A6C0;	14'h25B1: data <= 32'hE3EC381F;	14'h25B2: data <= 32'hE3F061B9;	14'h25B3: data <= 32'hE3F48B52;	14'h25B4: data <= 32'hE3F8B4EC;	14'h25B5: data <= 32'hE3FCDE86;	14'h25B6: data <= 32'hE401081F;	14'h25B7: data <= 32'hE40531B9;	14'h25B8: data <= 32'hE4095B53;	14'h25B9: data <= 32'hE40D84EC;	14'h25BA: data <= 32'hE411AE86;	14'h25BB: data <= 32'hE415D820;	14'h25BC: data <= 32'hE41A01B9;	14'h25BD: data <= 32'hE41E2B53;	14'h25BE: data <= 32'hE42254ED;	14'h25BF: data <= 32'hE4267E86;	14'h25C0: data <= 32'hE42AA820;	14'h25C1: data <= 32'hE42F287B;	14'h25C2: data <= 32'hE435D412;	14'h25C3: data <= 32'hE43C7FA9;	14'h25C4: data <= 32'hE4432B40;	14'h25C5: data <= 32'hE449D6D7;	14'h25C6: data <= 32'hE450826E;	14'h25C7: data <= 32'hE4572E05;	14'h25C8: data <= 32'hE45DD99C;	14'h25C9: data <= 32'hE4648533;	14'h25CA: data <= 32'hE46B30CA;	14'h25CB: data <= 32'hE471DC61;	14'h25CC: data <= 32'hE47887F8;	14'h25CD: data <= 32'hE47F338F;	14'h25CE: data <= 32'hE485DF26;	14'h25CF: data <= 32'hE48C8ABD;	14'h25D0: data <= 32'hE4933654;	14'h25D1: data <= 32'hE499E1EB;	14'h25D2: data <= 32'hE49C9360;	14'h25D3: data <= 32'hE49EEAFF;	14'h25D4: data <= 32'hE4A1429E;	14'h25D5: data <= 32'hE4A39A3C;	14'h25D6: data <= 32'hE4A5F1DB;	14'h25D7: data <= 32'hE4A8497A;	14'h25D8: data <= 32'hE4AAA119;	14'h25D9: data <= 32'hE4ACF8B7;	14'h25DA: data <= 32'hE4AF5056;	14'h25DB: data <= 32'hE4B1A7F5;	14'h25DC: data <= 32'hE4B3FF94;	14'h25DD: data <= 32'hE4B65732;	14'h25DE: data <= 32'hE4B8AED1;	14'h25DF: data <= 32'hE4BB0670;	14'h25E0: data <= 32'hE4BD5E0F;	14'h25E1: data <= 32'hE4BFB5AE;	14'h25E2: data <= 32'hE4BFCF08;	14'h25E3: data <= 32'hE4BEF56D;	14'h25E4: data <= 32'hE4BE1BD1;	14'h25E5: data <= 32'hE4BD4236;	14'h25E6: data <= 32'hE4BC689B;	14'h25E7: data <= 32'hE4BB8F00;	14'h25E8: data <= 32'hE4BAB565;	14'h25E9: data <= 32'hE4B9DBC9;	14'h25EA: data <= 32'hE4B9022E;	14'h25EB: data <= 32'hE4B82893;	14'h25EC: data <= 32'hE4B74EF8;	14'h25ED: data <= 32'hE4B6755D;	14'h25EE: data <= 32'hE4B59BC1;	14'h25EF: data <= 32'hE4B4C226;	14'h25F0: data <= 32'hE4B3E88B;	14'h25F1: data <= 32'hE4B30EF0;	14'h25F2: data <= 32'hE4B2E852;	14'h25F3: data <= 32'hE4B37EA2;	14'h25F4: data <= 32'hE4B414F2;	14'h25F5: data <= 32'hE4B4AB42;	14'h25F6: data <= 32'hE4B54193;	14'h25F7: data <= 32'hE4B5D7E3;	14'h25F8: data <= 32'hE4B66E33;	14'h25F9: data <= 32'hE4B70483;	14'h25FA: data <= 32'hE4B79AD4;	14'h25FB: data <= 32'hE4B83124;	14'h25FC: data <= 32'hE4B8C774;	14'h25FD: data <= 32'hE4B95DC4;	14'h25FE: data <= 32'hE4B9F415;	14'h25FF: data <= 32'hE4BA8A65;	14'h2600: data <= 32'hE4BB20B5;	14'h2601: data <= 32'hE4BBB705;	14'h2602: data <= 32'hE4BC721B;	14'h2603: data <= 32'hE4BD9077;	14'h2604: data <= 32'hE4BEAED3;	14'h2605: data <= 32'hE4BFCD2F;	14'h2606: data <= 32'hE4C0EB8B;	14'h2607: data <= 32'hE4C209E7;	14'h2608: data <= 32'hE4C32843;	14'h2609: data <= 32'hE4C446A0;	14'h260A: data <= 32'hE4C564FC;	14'h260B: data <= 32'hE4C68358;	14'h260C: data <= 32'hE4C7A1B4;	14'h260D: data <= 32'hE4C8C010;	14'h260E: data <= 32'hE4C9DE6C;	14'h260F: data <= 32'hE4CAFCC9;	14'h2610: data <= 32'hE4CC1B25;	14'h2611: data <= 32'hE4CD3981;	14'h2612: data <= 32'hE4CE76D9;	14'h2613: data <= 32'hE4D1D272;	14'h2614: data <= 32'hE4D52E0B;	14'h2615: data <= 32'hE4D889A3;	14'h2616: data <= 32'hE4DBE53C;	14'h2617: data <= 32'hE4DF40D5;	14'h2618: data <= 32'hE4E29C6D;	14'h2619: data <= 32'hE4E5F806;	14'h261A: data <= 32'hE4E9539F;	14'h261B: data <= 32'hE4ECAF37;	14'h261C: data <= 32'hE4F00AD0;	14'h261D: data <= 32'hE4F36668;	14'h261E: data <= 32'hE4F6C201;	14'h261F: data <= 32'hE4FA1D9A;	14'h2620: data <= 32'hE4FD7932;	14'h2621: data <= 32'hE500D4CB;	14'h2622: data <= 32'hE5043064;	14'h2623: data <= 32'hE5067182;	14'h2624: data <= 32'hE5087BF3;	14'h2625: data <= 32'hE50A8665;	14'h2626: data <= 32'hE50C90D7;	14'h2627: data <= 32'hE50E9B48;	14'h2628: data <= 32'hE510A5BA;	14'h2629: data <= 32'hE512B02B;	14'h262A: data <= 32'hE514BA9D;	14'h262B: data <= 32'hE516C50F;	14'h262C: data <= 32'hE518CF80;	14'h262D: data <= 32'hE51AD9F2;	14'h262E: data <= 32'hE51CE464;	14'h262F: data <= 32'hE51EEED5;	14'h2630: data <= 32'hE520F947;	14'h2631: data <= 32'hE52303B8;	14'h2632: data <= 32'hE5250E2A;	14'h2633: data <= 32'hE523921F;	14'h2634: data <= 32'hE51FF0BE;	14'h2635: data <= 32'hE51C4F5C;	14'h2636: data <= 32'hE518ADFB;	14'h2637: data <= 32'hE5150C99;	14'h2638: data <= 32'hE5116B37;	14'h2639: data <= 32'hE50DC9D6;	14'h263A: data <= 32'hE50A2874;	14'h263B: data <= 32'hE5068713;	14'h263C: data <= 32'hE502E5B1;	14'h263D: data <= 32'hE4FF444F;	14'h263E: data <= 32'hE4FBA2EE;	14'h263F: data <= 32'hE4F8018C;	14'h2640: data <= 32'hE4F4602B;	14'h2641: data <= 32'hE4F0BEC9;	14'h2642: data <= 32'hE4ED1D67;	14'h2643: data <= 32'hE4E85B1E;	14'h2644: data <= 32'hE4E1F11A;	14'h2645: data <= 32'hE4DB8716;	14'h2646: data <= 32'hE4D51D12;	14'h2647: data <= 32'hE4CEB30E;	14'h2648: data <= 32'hE4C84909;	14'h2649: data <= 32'hE4C1DF05;	14'h264A: data <= 32'hE4BB7501;	14'h264B: data <= 32'hE4B50AFD;	14'h264C: data <= 32'hE4AEA0F9;	14'h264D: data <= 32'hE4A836F5;	14'h264E: data <= 32'hE4A1CCF1;	14'h264F: data <= 32'hE49B62ED;	14'h2650: data <= 32'hE494F8E9;	14'h2651: data <= 32'hE48E8EE5;	14'h2652: data <= 32'hE48824E1;	14'h2653: data <= 32'hE481061F;	14'h2654: data <= 32'hE476E0C5;	14'h2655: data <= 32'hE46CBB6B;	14'h2656: data <= 32'hE4629611;	14'h2657: data <= 32'hE45870B7;	14'h2658: data <= 32'hE44E4B5D;	14'h2659: data <= 32'hE4442603;	14'h265A: data <= 32'hE43A00A9;	14'h265B: data <= 32'hE42FDB4E;	14'h265C: data <= 32'hE425B5F4;	14'h265D: data <= 32'hE41B909A;	14'h265E: data <= 32'hE4116B40;	14'h265F: data <= 32'hE40745E6;	14'h2660: data <= 32'hE3FD208C;	14'h2661: data <= 32'hE3F2FB32;	14'h2662: data <= 32'hE3E8D5D7;	14'h2663: data <= 32'hE3DEB07D;	14'h2664: data <= 32'hE3D79B3D;	14'h2665: data <= 32'hE3D09BC5;	14'h2666: data <= 32'hE3C99C4D;	14'h2667: data <= 32'hE3C29CD5;	14'h2668: data <= 32'hE3BB9D5C;	14'h2669: data <= 32'hE3B49DE4;	14'h266A: data <= 32'hE3AD9E6C;	14'h266B: data <= 32'hE3A69EF4;	14'h266C: data <= 32'hE39F9F7B;	14'h266D: data <= 32'hE398A003;	14'h266E: data <= 32'hE391A08B;	14'h266F: data <= 32'hE38AA113;	14'h2670: data <= 32'hE383A19A;	14'h2671: data <= 32'hE37CA222;	14'h2672: data <= 32'hE375A2AA;	14'h2673: data <= 32'hE36EA332;	14'h2674: data <= 32'hE369D298;	14'h2675: data <= 32'hE365B5A0;	14'h2676: data <= 32'hE36198A9;	14'h2677: data <= 32'hE35D7BB1;	14'h2678: data <= 32'hE3595EBA;	14'h2679: data <= 32'hE35541C2;	14'h267A: data <= 32'hE35124CB;	14'h267B: data <= 32'hE34D07D4;	14'h267C: data <= 32'hE348EADC;	14'h267D: data <= 32'hE344CDE5;	14'h267E: data <= 32'hE340B0ED;	14'h267F: data <= 32'hE33C93F6;	14'h2680: data <= 32'hE33876FE;	14'h2681: data <= 32'hE3345A07;	14'h2682: data <= 32'hE3303D10;	14'h2683: data <= 32'hE32C2018;	14'h2684: data <= 32'hE32762FF;	14'h2685: data <= 32'hE3221DC9;	14'h2686: data <= 32'hE31CD893;	14'h2687: data <= 32'hE317935E;	14'h2688: data <= 32'hE3124E28;	14'h2689: data <= 32'hE30D08F2;	14'h268A: data <= 32'hE307C3BC;	14'h268B: data <= 32'hE3027E87;	14'h268C: data <= 32'hE2FD3951;	14'h268D: data <= 32'hE2F7F41B;	14'h268E: data <= 32'hE2F2AEE5;	14'h268F: data <= 32'hE2ED69AF;	14'h2690: data <= 32'hE2E8247A;	14'h2691: data <= 32'hE2E2DF44;	14'h2692: data <= 32'hE2DD9A0E;	14'h2693: data <= 32'hE2D854D8;	14'h2694: data <= 32'hE2D46A21;	14'h2695: data <= 32'hE2D35144;	14'h2696: data <= 32'hE2D23868;	14'h2697: data <= 32'hE2D11F8C;	14'h2698: data <= 32'hE2D006B0;	14'h2699: data <= 32'hE2CEEDD4;	14'h269A: data <= 32'hE2CDD4F8;	14'h269B: data <= 32'hE2CCBC1C;	14'h269C: data <= 32'hE2CBA340;	14'h269D: data <= 32'hE2CA8A63;	14'h269E: data <= 32'hE2C97187;	14'h269F: data <= 32'hE2C858AB;	14'h26A0: data <= 32'hE2C73FCF;	14'h26A1: data <= 32'hE2C626F3;	14'h26A2: data <= 32'hE2C50E17;	14'h26A3: data <= 32'hE2C3F53B;	14'h26A4: data <= 32'hE2C3172C;	14'h26A5: data <= 32'hE2C41E3E;	14'h26A6: data <= 32'hE2C52550;	14'h26A7: data <= 32'hE2C62C62;	14'h26A8: data <= 32'hE2C73374;	14'h26A9: data <= 32'hE2C83A85;	14'h26AA: data <= 32'hE2C94197;	14'h26AB: data <= 32'hE2CA48A9;	14'h26AC: data <= 32'hE2CB4FBB;	14'h26AD: data <= 32'hE2CC56CD;	14'h26AE: data <= 32'hE2CD5DDF;	14'h26AF: data <= 32'hE2CE64F1;	14'h26B0: data <= 32'hE2CF6C02;	14'h26B1: data <= 32'hE2D07314;	14'h26B2: data <= 32'hE2D17A26;	14'h26B3: data <= 32'hE2D28138;	14'h26B4: data <= 32'hE2D3884A;	14'h26B5: data <= 32'hE2D5BFAA;	14'h26B6: data <= 32'hE2D81BED;	14'h26B7: data <= 32'hE2DA7830;	14'h26B8: data <= 32'hE2DCD472;	14'h26B9: data <= 32'hE2DF30B5;	14'h26BA: data <= 32'hE2E18CF8;	14'h26BB: data <= 32'hE2E3E93B;	14'h26BC: data <= 32'hE2E6457E;	14'h26BD: data <= 32'hE2E8A1C1;	14'h26BE: data <= 32'hE2EAFE03;	14'h26BF: data <= 32'hE2ED5A46;	14'h26C0: data <= 32'hE2EFB689;	14'h26C1: data <= 32'hE2F212CC;	14'h26C2: data <= 32'hE2F46F0F;	14'h26C3: data <= 32'hE2F6CB52;	14'h26C4: data <= 32'hE2F92794;	14'h26C5: data <= 32'hE2FEB1EA;	14'h26C6: data <= 32'hE305C300;	14'h26C7: data <= 32'hE30CD417;	14'h26C8: data <= 32'hE313E52D;	14'h26C9: data <= 32'hE31AF644;	14'h26CA: data <= 32'hE322075A;	14'h26CB: data <= 32'hE3291871;	14'h26CC: data <= 32'hE3302988;	14'h26CD: data <= 32'hE3373A9E;	14'h26CE: data <= 32'hE33E4BB5;	14'h26CF: data <= 32'hE3455CCB;	14'h26D0: data <= 32'hE34C6DE2;	14'h26D1: data <= 32'hE3537EF8;	14'h26D2: data <= 32'hE35A900F;	14'h26D3: data <= 32'hE361A125;	14'h26D4: data <= 32'hE368B23C;	14'h26D5: data <= 32'hE37245E5;	14'h26D6: data <= 32'hE37ECD86;	14'h26D7: data <= 32'hE38B5527;	14'h26D8: data <= 32'hE397DCC8;	14'h26D9: data <= 32'hE3A46469;	14'h26DA: data <= 32'hE3B0EC0A;	14'h26DB: data <= 32'hE3BD73AB;	14'h26DC: data <= 32'hE3C9FB4C;	14'h26DD: data <= 32'hE3D682ED;	14'h26DE: data <= 32'hE3E30A8E;	14'h26DF: data <= 32'hE3EF922F;	14'h26E0: data <= 32'hE3FC19D0;	14'h26E1: data <= 32'hE408A171;	14'h26E2: data <= 32'hE4152912;	14'h26E3: data <= 32'hE421B0B3;	14'h26E4: data <= 32'hE42E3854;	14'h26E5: data <= 32'hE43B6E2E;	14'h26E6: data <= 32'hE44AC20E;	14'h26E7: data <= 32'hE45A15ED;	14'h26E8: data <= 32'hE46969CD;	14'h26E9: data <= 32'hE478BDAC;	14'h26EA: data <= 32'hE488118C;	14'h26EB: data <= 32'hE497656B;	14'h26EC: data <= 32'hE4A6B94B;	14'h26ED: data <= 32'hE4B60D2A;	14'h26EE: data <= 32'hE4C5610A;	14'h26EF: data <= 32'hE4D4B4E9;	14'h26F0: data <= 32'hE4E408C9;	14'h26F1: data <= 32'hE4F35CA8;	14'h26F2: data <= 32'hE502B088;	14'h26F3: data <= 32'hE5120467;	14'h26F4: data <= 32'hE5215847;	14'h26F5: data <= 32'hE530AA2C;	14'h26F6: data <= 32'hE53FB4E9;	14'h26F7: data <= 32'hE54EBFA5;	14'h26F8: data <= 32'hE55DCA62;	14'h26F9: data <= 32'hE56CD51E;	14'h26FA: data <= 32'hE57BDFDB;	14'h26FB: data <= 32'hE58AEA97;	14'h26FC: data <= 32'hE599F554;	14'h26FD: data <= 32'hE5A90010;	14'h26FE: data <= 32'hE5B80ACD;	14'h26FF: data <= 32'hE5C71589;	14'h2700: data <= 32'hE5D62046;	14'h2701: data <= 32'hE5E52B02;	14'h2702: data <= 32'hE5F435BF;	14'h2703: data <= 32'hE603407B;	14'h2704: data <= 32'hE6124B38;	14'h2705: data <= 32'hE62155F4;	14'h2706: data <= 32'hE62B7431;	14'h2707: data <= 32'hE6346C51;	14'h2708: data <= 32'hE63D6471;	14'h2709: data <= 32'hE6465C90;	14'h270A: data <= 32'hE64F54B0;	14'h270B: data <= 32'hE6584CD0;	14'h270C: data <= 32'hE66144EF;	14'h270D: data <= 32'hE66A3D0F;	14'h270E: data <= 32'hE673352F;	14'h270F: data <= 32'hE67C2D4E;	14'h2710: data <= 32'hE685256E;	14'h2711: data <= 32'hE68E1D8D;	14'h2712: data <= 32'hE69715AD;	14'h2713: data <= 32'hE6A00DCD;	14'h2714: data <= 32'hE6A905EC;	14'h2715: data <= 32'hE6B1FE0C;	14'h2716: data <= 32'hE6B7288C;	14'h2717: data <= 32'hE6B9BB35;	14'h2718: data <= 32'hE6BC4DDF;	14'h2719: data <= 32'hE6BEE089;	14'h271A: data <= 32'hE6C17332;	14'h271B: data <= 32'hE6C405DC;	14'h271C: data <= 32'hE6C69886;	14'h271D: data <= 32'hE6C92B30;	14'h271E: data <= 32'hE6CBBDD9;	14'h271F: data <= 32'hE6CE5083;	14'h2720: data <= 32'hE6D0E32D;	14'h2721: data <= 32'hE6D375D6;	14'h2722: data <= 32'hE6D60880;	14'h2723: data <= 32'hE6D89B2A;	14'h2724: data <= 32'hE6DB2DD3;	14'h2725: data <= 32'hE6DDC07D;	14'h2726: data <= 32'hE6DE0511;	14'h2727: data <= 32'hE6DA8038;	14'h2728: data <= 32'hE6D6FB5E;	14'h2729: data <= 32'hE6D37685;	14'h272A: data <= 32'hE6CFF1AC;	14'h272B: data <= 32'hE6CC6CD3;	14'h272C: data <= 32'hE6C8E7F9;	14'h272D: data <= 32'hE6C56320;	14'h272E: data <= 32'hE6C1DE47;	14'h272F: data <= 32'hE6BE596E;	14'h2730: data <= 32'hE6BAD495;	14'h2731: data <= 32'hE6B74FBB;	14'h2732: data <= 32'hE6B3CAE2;	14'h2733: data <= 32'hE6B04609;	14'h2734: data <= 32'hE6ACC130;	14'h2735: data <= 32'hE6A93C56;	14'h2736: data <= 32'hE6A53725;	14'h2737: data <= 32'hE69E9ADB;	14'h2738: data <= 32'hE697FE90;	14'h2739: data <= 32'hE6916245;	14'h273A: data <= 32'hE68AC5FA;	14'h273B: data <= 32'hE68429AF;	14'h273C: data <= 32'hE67D8D64;	14'h273D: data <= 32'hE676F11A;	14'h273E: data <= 32'hE67054CF;	14'h273F: data <= 32'hE669B884;	14'h2740: data <= 32'hE6631C39;	14'h2741: data <= 32'hE65C7FEE;	14'h2742: data <= 32'hE655E3A3;	14'h2743: data <= 32'hE64F4759;	14'h2744: data <= 32'hE648AB0E;	14'h2745: data <= 32'hE6420EC3;	14'h2746: data <= 32'hE63B7278;	14'h2747: data <= 32'hE63796C7;	14'h2748: data <= 32'hE633E359;	14'h2749: data <= 32'hE6302FEB;	14'h274A: data <= 32'hE62C7C7D;	14'h274B: data <= 32'hE628C910;	14'h274C: data <= 32'hE62515A2;	14'h274D: data <= 32'hE6216234;	14'h274E: data <= 32'hE61DAEC6;	14'h274F: data <= 32'hE619FB58;	14'h2750: data <= 32'hE61647EA;	14'h2751: data <= 32'hE612947D;	14'h2752: data <= 32'hE60EE10F;	14'h2753: data <= 32'hE60B2DA1;	14'h2754: data <= 32'hE6077A33;	14'h2755: data <= 32'hE603C6C5;	14'h2756: data <= 32'hE6001357;	14'h2757: data <= 32'hE5FF35E6;	14'h2758: data <= 32'hE5FF6557;	14'h2759: data <= 32'hE5FF94C7;	14'h275A: data <= 32'hE5FFC438;	14'h275B: data <= 32'hE5FFF3A9;	14'h275C: data <= 32'hE6002319;	14'h275D: data <= 32'hE600528A;	14'h275E: data <= 32'hE60081FB;	14'h275F: data <= 32'hE600B16B;	14'h2760: data <= 32'hE600E0DC;	14'h2761: data <= 32'hE601104D;	14'h2762: data <= 32'hE6013FBD;	14'h2763: data <= 32'hE6016F2E;	14'h2764: data <= 32'hE6019E9F;	14'h2765: data <= 32'hE601CE10;	14'h2766: data <= 32'hE601FD80;	14'h2767: data <= 32'hE60222E1;	14'h2768: data <= 32'hE6023EB9;	14'h2769: data <= 32'hE6025A92;	14'h276A: data <= 32'hE602766A;	14'h276B: data <= 32'hE6029243;	14'h276C: data <= 32'hE602AE1B;	14'h276D: data <= 32'hE602C9F4;	14'h276E: data <= 32'hE602E5CC;	14'h276F: data <= 32'hE60301A4;	14'h2770: data <= 32'hE6031D7D;	14'h2771: data <= 32'hE6033955;	14'h2772: data <= 32'hE603552E;	14'h2773: data <= 32'hE6037106;	14'h2774: data <= 32'hE6038CDE;	14'h2775: data <= 32'hE603A8B7;	14'h2776: data <= 32'hE603C48F;	14'h2777: data <= 32'hE60319C7;	14'h2778: data <= 32'hE6009981;	14'h2779: data <= 32'hE5FE193C;	14'h277A: data <= 32'hE5FB98F7;	14'h277B: data <= 32'hE5F918B1;	14'h277C: data <= 32'hE5F6986C;	14'h277D: data <= 32'hE5F41826;	14'h277E: data <= 32'hE5F197E1;	14'h277F: data <= 32'hE5EF179C;	14'h2780: data <= 32'hE5EC9756;	14'h2781: data <= 32'hE5EA1711;	14'h2782: data <= 32'hE5E796CB;	14'h2783: data <= 32'hE5E51686;	14'h2784: data <= 32'hE5E29641;	14'h2785: data <= 32'hE5E015FB;	14'h2786: data <= 32'hE5DD95B6;	14'h2787: data <= 32'hE5DAC4E3;	14'h2788: data <= 32'hE5D4631F;	14'h2789: data <= 32'hE5CE015B;	14'h278A: data <= 32'hE5C79F97;	14'h278B: data <= 32'hE5C13DD3;	14'h278C: data <= 32'hE5BADC0F;	14'h278D: data <= 32'hE5B47A4B;	14'h278E: data <= 32'hE5AE1887;	14'h278F: data <= 32'hE5A7B6C3;	14'h2790: data <= 32'hE5A154FF;	14'h2791: data <= 32'hE59AF33B;	14'h2792: data <= 32'hE5949177;	14'h2793: data <= 32'hE58E2FB3;	14'h2794: data <= 32'hE587CDEF;	14'h2795: data <= 32'hE5816C2B;	14'h2796: data <= 32'hE57B0A67;	14'h2797: data <= 32'hE574A8A3;	14'h2798: data <= 32'hE56C9387;	14'h2799: data <= 32'hE5643A66;	14'h279A: data <= 32'hE55BE145;	14'h279B: data <= 32'hE5538823;	14'h279C: data <= 32'hE54B2F02;	14'h279D: data <= 32'hE542D5E1;	14'h279E: data <= 32'hE53A7CBF;	14'h279F: data <= 32'hE532239E;	14'h27A0: data <= 32'hE529CA7D;	14'h27A1: data <= 32'hE521715C;	14'h27A2: data <= 32'hE519183A;	14'h27A3: data <= 32'hE510BF19;	14'h27A4: data <= 32'hE50865F8;	14'h27A5: data <= 32'hE5000CD6;	14'h27A6: data <= 32'hE4F7B3B5;	14'h27A7: data <= 32'hE4EF5A94;	14'h27A8: data <= 32'hE4E6C1F4;	14'h27A9: data <= 32'hE4DE06EF;	14'h27AA: data <= 32'hE4D54BEA;	14'h27AB: data <= 32'hE4CC90E5;	14'h27AC: data <= 32'hE4C3D5E0;	14'h27AD: data <= 32'hE4BB1ADC;	14'h27AE: data <= 32'hE4B25FD7;	14'h27AF: data <= 32'hE4A9A4D2;	14'h27B0: data <= 32'hE4A0E9CD;	14'h27B1: data <= 32'hE4982EC8;	14'h27B2: data <= 32'hE48F73C4;	14'h27B3: data <= 32'hE486B8BF;	14'h27B4: data <= 32'hE47DFDBA;	14'h27B5: data <= 32'hE47542B5;	14'h27B6: data <= 32'hE46C87B0;	14'h27B7: data <= 32'hE463CCAC;	14'h27B8: data <= 32'hE45C3421;	14'h27B9: data <= 32'hE45618D6;	14'h27BA: data <= 32'hE44FFD8B;	14'h27BB: data <= 32'hE449E240;	14'h27BC: data <= 32'hE443C6F5;	14'h27BD: data <= 32'hE43DABAA;	14'h27BE: data <= 32'hE437905F;	14'h27BF: data <= 32'hE4317514;	14'h27C0: data <= 32'hE42B59C9;	14'h27C1: data <= 32'hE4253E7F;	14'h27C2: data <= 32'hE41F2334;	14'h27C3: data <= 32'hE41907E9;	14'h27C4: data <= 32'hE412EC9E;	14'h27C5: data <= 32'hE40CD153;	14'h27C6: data <= 32'hE406B608;	14'h27C7: data <= 32'hE4009ABD;	14'h27C8: data <= 32'hE3FB196B;	14'h27C9: data <= 32'hE3F7C63E;	14'h27CA: data <= 32'hE3F47312;	14'h27CB: data <= 32'hE3F11FE6;	14'h27CC: data <= 32'hE3EDCCB9;	14'h27CD: data <= 32'hE3EA798D;	14'h27CE: data <= 32'hE3E72660;	14'h27CF: data <= 32'hE3E3D334;	14'h27D0: data <= 32'hE3E08007;	14'h27D1: data <= 32'hE3DD2CDB;	14'h27D2: data <= 32'hE3D9D9AE;	14'h27D3: data <= 32'hE3D68682;	14'h27D4: data <= 32'hE3D33355;	14'h27D5: data <= 32'hE3CFE029;	14'h27D6: data <= 32'hE3CC8CFC;	14'h27D7: data <= 32'hE3C939D0;	14'h27D8: data <= 32'hE3C5E6A3;	14'h27D9: data <= 32'hE3C312EB;	14'h27DA: data <= 32'hE3C03F32;	14'h27DB: data <= 32'hE3BD6B7A;	14'h27DC: data <= 32'hE3BA97C1;	14'h27DD: data <= 32'hE3B7C408;	14'h27DE: data <= 32'hE3B4F050;	14'h27DF: data <= 32'hE3B21C97;	14'h27E0: data <= 32'hE3AF48DE;	14'h27E1: data <= 32'hE3AC7526;	14'h27E2: data <= 32'hE3A9A16D;	14'h27E3: data <= 32'hE3A6CDB5;	14'h27E4: data <= 32'hE3A3F9FC;	14'h27E5: data <= 32'hE3A12643;	14'h27E6: data <= 32'hE39E528B;	14'h27E7: data <= 32'hE39B7ED2;	14'h27E8: data <= 32'hE398AB19;	14'h27E9: data <= 32'hE3947589;	14'h27EA: data <= 32'hE38FDE5C;	14'h27EB: data <= 32'hE38B472E;	14'h27EC: data <= 32'hE386B001;	14'h27ED: data <= 32'hE38218D4;	14'h27EE: data <= 32'hE37D81A7;	14'h27EF: data <= 32'hE378EA7A;	14'h27F0: data <= 32'hE374534C;	14'h27F1: data <= 32'hE36FBC1F;	14'h27F2: data <= 32'hE36B24F2;	14'h27F3: data <= 32'hE3668DC5;	14'h27F4: data <= 32'hE361F698;	14'h27F5: data <= 32'hE35D5F6A;	14'h27F6: data <= 32'hE358C83D;	14'h27F7: data <= 32'hE3543110;	14'h27F8: data <= 32'hE34F99E3;	14'h27F9: data <= 32'hE34C5379;	14'h27FA: data <= 32'hE34A0DA5;	14'h27FB: data <= 32'hE347C7D0;	14'h27FC: data <= 32'hE34581FB;	14'h27FD: data <= 32'hE3433C27;	14'h27FE: data <= 32'hE340F652;	14'h27FF: data <= 32'hE33EB07E;	14'h2800: data <= 32'hE33C6AA9;	14'h2801: data <= 32'hE33A24D5;	14'h2802: data <= 32'hE337DF00;	14'h2803: data <= 32'hE335992C;	14'h2804: data <= 32'hE3335357;	14'h2805: data <= 32'hE3310D82;	14'h2806: data <= 32'hE32EC7AE;	14'h2807: data <= 32'hE32C81D9;	14'h2808: data <= 32'hE32A3C05;	14'h2809: data <= 32'hE3291CDF;	14'h280A: data <= 32'hE32A1DC1;	14'h280B: data <= 32'hE32B1EA3;	14'h280C: data <= 32'hE32C1F84;	14'h280D: data <= 32'hE32D2066;	14'h280E: data <= 32'hE32E2148;	14'h280F: data <= 32'hE32F222A;	14'h2810: data <= 32'hE330230B;	14'h2811: data <= 32'hE33123ED;	14'h2812: data <= 32'hE33224CF;	14'h2813: data <= 32'hE33325B1;	14'h2814: data <= 32'hE3342692;	14'h2815: data <= 32'hE3352774;	14'h2816: data <= 32'hE3362856;	14'h2817: data <= 32'hE3372938;	14'h2818: data <= 32'hE3382A19;	14'h2819: data <= 32'hE3393821;	14'h281A: data <= 32'hE33A9A4C;	14'h281B: data <= 32'hE33BFC77;	14'h281C: data <= 32'hE33D5EA2;	14'h281D: data <= 32'hE33EC0CE;	14'h281E: data <= 32'hE34022F9;	14'h281F: data <= 32'hE3418524;	14'h2820: data <= 32'hE342E74F;	14'h2821: data <= 32'hE344497A;	14'h2822: data <= 32'hE345ABA6;	14'h2823: data <= 32'hE3470DD1;	14'h2824: data <= 32'hE3486FFC;	14'h2825: data <= 32'hE349D227;	14'h2826: data <= 32'hE34B3452;	14'h2827: data <= 32'hE34C967E;	14'h2828: data <= 32'hE34DF8A9;	14'h2829: data <= 32'hE34F5AD4;	14'h282A: data <= 32'hE34E11F3;	14'h282B: data <= 32'hE34C8CCE;	14'h282C: data <= 32'hE34B07A8;	14'h282D: data <= 32'hE3498282;	14'h282E: data <= 32'hE347FD5C;	14'h282F: data <= 32'hE3467837;	14'h2830: data <= 32'hE344F311;	14'h2831: data <= 32'hE3436DEB;	14'h2832: data <= 32'hE341E8C6;	14'h2833: data <= 32'hE34063A0;	14'h2834: data <= 32'hE33EDE7A;	14'h2835: data <= 32'hE33D5955;	14'h2836: data <= 32'hE33BD42F;	14'h2837: data <= 32'hE33A4F09;	14'h2838: data <= 32'hE338C9E3;	14'h2839: data <= 32'hE33744BE;	14'h283A: data <= 32'hE32F2D9E;	14'h283B: data <= 32'hE3244EE3;	14'h283C: data <= 32'hE3197028;	14'h283D: data <= 32'hE30E916E;	14'h283E: data <= 32'hE303B2B3;	14'h283F: data <= 32'hE2F8D3F8;	14'h2840: data <= 32'hE2EDF53D;	14'h2841: data <= 32'hE2E31682;	14'h2842: data <= 32'hE2D837C7;	14'h2843: data <= 32'hE2CD590D;	14'h2844: data <= 32'hE2C27A52;	14'h2845: data <= 32'hE2B79B97;	14'h2846: data <= 32'hE2ACBCDC;	14'h2847: data <= 32'hE2A1DE21;	14'h2848: data <= 32'hE296FF66;	14'h2849: data <= 32'hE28C20AC;	14'h284A: data <= 32'hE27FFA3C;	14'h284B: data <= 32'hE27279E4;	14'h284C: data <= 32'hE264F98B;	14'h284D: data <= 32'hE2577932;	14'h284E: data <= 32'hE249F8DA;	14'h284F: data <= 32'hE23C7881;	14'h2850: data <= 32'hE22EF828;	14'h2851: data <= 32'hE22177D0;	14'h2852: data <= 32'hE213F777;	14'h2853: data <= 32'hE206771E;	14'h2854: data <= 32'hE1F8F6C6;	14'h2855: data <= 32'hE1EB766D;	14'h2856: data <= 32'hE1DDF614;	14'h2857: data <= 32'hE1D075BC;	14'h2858: data <= 32'hE1C2F563;	14'h2859: data <= 32'hE1B5750A;	14'h285A: data <= 32'hE1A76EBD;	14'h285B: data <= 32'hE197FEC4;	14'h285C: data <= 32'hE1888ECA;	14'h285D: data <= 32'hE1791ED0;	14'h285E: data <= 32'hE169AED6;	14'h285F: data <= 32'hE15A3EDC;	14'h2860: data <= 32'hE14ACEE2;	14'h2861: data <= 32'hE13B5EE8;	14'h2862: data <= 32'hE12BEEEE;	14'h2863: data <= 32'hE11C7EF4;	14'h2864: data <= 32'hE10D0EFA;	14'h2865: data <= 32'hE0FD9F00;	14'h2866: data <= 32'hE0EE2F06;	14'h2867: data <= 32'hE0DEBF0C;	14'h2868: data <= 32'hE0CF4F13;	14'h2869: data <= 32'hE0BFDF19;	14'h286A: data <= 32'hE0AFB9DD;	14'h286B: data <= 32'hE09330AC;	14'h286C: data <= 32'hE076A77B;	14'h286D: data <= 32'hE05A1E4A;	14'h286E: data <= 32'hE03D9519;	14'h286F: data <= 32'hE0210BE8;	14'h2870: data <= 32'hE00482B7;	14'h2871: data <= 32'hDFE7F986;	14'h2872: data <= 32'hDFCB7055;	14'h2873: data <= 32'hDFAEE723;	14'h2874: data <= 32'hDF925DF2;	14'h2875: data <= 32'hDF75D4C1;	14'h2876: data <= 32'hDF594B90;	14'h2877: data <= 32'hDF3CC25F;	14'h2878: data <= 32'hDF20392E;	14'h2879: data <= 32'hDF03AFFD;	14'h287A: data <= 32'hDEE726CC;	14'h287B: data <= 32'hDEC28107;	14'h287C: data <= 32'hDE9C4958;	14'h287D: data <= 32'hDE7611A8;	14'h287E: data <= 32'hDE4FD9F9;	14'h287F: data <= 32'hDE29A24A;	14'h2880: data <= 32'hDE036A9A;	14'h2881: data <= 32'hDDDD32EB;	14'h2882: data <= 32'hDDB6FB3B;	14'h2883: data <= 32'hDD90C38C;	14'h2884: data <= 32'hDD6A8BDC;	14'h2885: data <= 32'hDD44542D;	14'h2886: data <= 32'hDD1E1C7E;	14'h2887: data <= 32'hDCF7E4CE;	14'h2888: data <= 32'hDCD1AD1F;	14'h2889: data <= 32'hDCAB756F;	14'h288A: data <= 32'hDC853DC0;	14'h288B: data <= 32'hDC63F819;	14'h288C: data <= 32'hDC45B514;	14'h288D: data <= 32'hDC27720E;	14'h288E: data <= 32'hDC092F08;	14'h288F: data <= 32'hDBEAEC03;	14'h2890: data <= 32'hDBCCA8FD;	14'h2891: data <= 32'hDBAE65F7;	14'h2892: data <= 32'hDB9022F2;	14'h2893: data <= 32'hDB71DFEC;	14'h2894: data <= 32'hDB539CE7;	14'h2895: data <= 32'hDB3559E1;	14'h2896: data <= 32'hDB1716DB;	14'h2897: data <= 32'hDAF8D3D6;	14'h2898: data <= 32'hDADA90D0;	14'h2899: data <= 32'hDABC4DCA;	14'h289A: data <= 32'hDA9E0AC5;	14'h289B: data <= 32'hDA8440C7;	14'h289C: data <= 32'hDA71062B;	14'h289D: data <= 32'hDA5DCB8F;	14'h289E: data <= 32'hDA4A90F3;	14'h289F: data <= 32'hDA375657;	14'h28A0: data <= 32'hDA241BBA;	14'h28A1: data <= 32'hDA10E11E;	14'h28A2: data <= 32'hD9FDA682;	14'h28A3: data <= 32'hD9EA6BE6;	14'h28A4: data <= 32'hD9D7314A;	14'h28A5: data <= 32'hD9C3F6AE;	14'h28A6: data <= 32'hD9B0BC11;	14'h28A7: data <= 32'hD99D8175;	14'h28A8: data <= 32'hD98A46D9;	14'h28A9: data <= 32'hD9770C3D;	14'h28AA: data <= 32'hD963D1A1;	14'h28AB: data <= 32'hD9521A1F;	14'h28AC: data <= 32'hD946DDA1;	14'h28AD: data <= 32'hD93BA123;	14'h28AE: data <= 32'hD93064A5;	14'h28AF: data <= 32'hD9252826;	14'h28B0: data <= 32'hD919EBA8;	14'h28B1: data <= 32'hD90EAF2A;	14'h28B2: data <= 32'hD90372AC;	14'h28B3: data <= 32'hD8F8362E;	14'h28B4: data <= 32'hD8ECF9B0;	14'h28B5: data <= 32'hD8E1BD32;	14'h28B6: data <= 32'hD8D680B3;	14'h28B7: data <= 32'hD8CB4435;	14'h28B8: data <= 32'hD8C007B7;	14'h28B9: data <= 32'hD8B4CB39;	14'h28BA: data <= 32'hD8A98EBB;	14'h28BB: data <= 32'hD89E523D;	14'h28BC: data <= 32'hD88C8B18;	14'h28BD: data <= 32'hD87A956F;	14'h28BE: data <= 32'hD8689FC5;	14'h28BF: data <= 32'hD856AA1C;	14'h28C0: data <= 32'hD844B472;	14'h28C1: data <= 32'hD832BEC9;	14'h28C2: data <= 32'hD820C920;	14'h28C3: data <= 32'hD80ED376;	14'h28C4: data <= 32'hD7FCDDCD;	14'h28C5: data <= 32'hD7EAE823;	14'h28C6: data <= 32'hD7D8F27A;	14'h28C7: data <= 32'hD7C6FCD1;	14'h28C8: data <= 32'hD7B50727;	14'h28C9: data <= 32'hD7A3117E;	14'h28CA: data <= 32'hD7911BD5;	14'h28CB: data <= 32'hD77F262B;	14'h28CC: data <= 32'hD75FBDD0;	14'h28CD: data <= 32'hD73C02DF;	14'h28CE: data <= 32'hD71847EF;	14'h28CF: data <= 32'hD6F48CFF;	14'h28D0: data <= 32'hD6D0D20F;	14'h28D1: data <= 32'hD6AD171F;	14'h28D2: data <= 32'hD6895C2F;	14'h28D3: data <= 32'hD665A13F;	14'h28D4: data <= 32'hD641E64E;	14'h28D5: data <= 32'hD61E2B5E;	14'h28D6: data <= 32'hD5FA706E;	14'h28D7: data <= 32'hD5D6B57E;	14'h28D8: data <= 32'hD5B2FA8E;	14'h28D9: data <= 32'hD58F3F9E;	14'h28DA: data <= 32'hD56B84AD;	14'h28DB: data <= 32'hD547C9BD;	14'h28DC: data <= 32'hD5207C18;	14'h28DD: data <= 32'hD4F624F3;	14'h28DE: data <= 32'hD4CBCDCF;	14'h28DF: data <= 32'hD4A176AA;	14'h28E0: data <= 32'hD4771F85;	14'h28E1: data <= 32'hD44CC860;	14'h28E2: data <= 32'hD422713B;	14'h28E3: data <= 32'hD3F81A16;	14'h28E4: data <= 32'hD3CDC2F1;	14'h28E5: data <= 32'hD3A36BCD;	14'h28E6: data <= 32'hD37914A8;	14'h28E7: data <= 32'hD34EBD83;	14'h28E8: data <= 32'hD324665E;	14'h28E9: data <= 32'hD2FA0F39;	14'h28EA: data <= 32'hD2CFB814;	14'h28EB: data <= 32'hD2A560EF;	14'h28EC: data <= 32'hD27FB571;	14'h28ED: data <= 32'hD263C4E2;	14'h28EE: data <= 32'hD247D453;	14'h28EF: data <= 32'hD22BE3C4;	14'h28F0: data <= 32'hD20FF335;	14'h28F1: data <= 32'hD1F402A6;	14'h28F2: data <= 32'hD1D81218;	14'h28F3: data <= 32'hD1BC2189;	14'h28F4: data <= 32'hD1A030FA;	14'h28F5: data <= 32'hD184406B;	14'h28F6: data <= 32'hD1684FDC;	14'h28F7: data <= 32'hD14C5F4D;	14'h28F8: data <= 32'hD1306EBE;	14'h28F9: data <= 32'hD1147E2F;	14'h28FA: data <= 32'hD0F88DA0;	14'h28FB: data <= 32'hD0DC9D12;	14'h28FC: data <= 32'hD0C1B362;	14'h28FD: data <= 32'hD0AF4265;	14'h28FE: data <= 32'hD09CD167;	14'h28FF: data <= 32'hD08A606A;	14'h2900: data <= 32'hD077EF6D;	14'h2901: data <= 32'hD0657E70;	14'h2902: data <= 32'hD0530D72;	14'h2903: data <= 32'hD0409C75;	14'h2904: data <= 32'hD02E2B78;	14'h2905: data <= 32'hD01BBA7B;	14'h2906: data <= 32'hD009497E;	14'h2907: data <= 32'hCFF6D880;	14'h2908: data <= 32'hCFE46783;	14'h2909: data <= 32'hCFD1F686;	14'h290A: data <= 32'hCFBF8589;	14'h290B: data <= 32'hCFAD148B;	14'h290C: data <= 32'hCF9AA38E;	14'h290D: data <= 32'hCF88E6ED;	14'h290E: data <= 32'hCF774029;	14'h290F: data <= 32'hCF659965;	14'h2910: data <= 32'hCF53F2A0;	14'h2911: data <= 32'hCF424BDC;	14'h2912: data <= 32'hCF30A518;	14'h2913: data <= 32'hCF1EFE54;	14'h2914: data <= 32'hCF0D578F;	14'h2915: data <= 32'hCEFBB0CB;	14'h2916: data <= 32'hCEEA0A07;	14'h2917: data <= 32'hCED86343;	14'h2918: data <= 32'hCEC6BC7E;	14'h2919: data <= 32'hCEB515BA;	14'h291A: data <= 32'hCEA36EF6;	14'h291B: data <= 32'hCE91C832;	14'h291C: data <= 32'hCE80216D;	14'h291D: data <= 32'hCE629FF7;	14'h291E: data <= 32'hCE3F6DD9;	14'h291F: data <= 32'hCE1C3BBB;	14'h2920: data <= 32'hCDF9099D;	14'h2921: data <= 32'hCDD5D77F;	14'h2922: data <= 32'hCDB2A560;	14'h2923: data <= 32'hCD8F7342;	14'h2924: data <= 32'hCD6C4124;	14'h2925: data <= 32'hCD490F06;	14'h2926: data <= 32'hCD25DCE8;	14'h2927: data <= 32'hCD02AACA;	14'h2928: data <= 32'hCCDF78AC;	14'h2929: data <= 32'hCCBC468E;	14'h292A: data <= 32'hCC991470;	14'h292B: data <= 32'hCC75E252;	14'h292C: data <= 32'hCC52B034;	14'h292D: data <= 32'hCC1A54A9;	14'h292E: data <= 32'hCBC913AC;	14'h292F: data <= 32'hCB77D2AE;	14'h2930: data <= 32'hCB2691B1;	14'h2931: data <= 32'hCAD550B4;	14'h2932: data <= 32'hCA840FB7;	14'h2933: data <= 32'hCA32CEBA;	14'h2934: data <= 32'hC9E18DBD;	14'h2935: data <= 32'hC9904CC0;	14'h2936: data <= 32'hC93F0BC3;	14'h2937: data <= 32'hC8EDCAC6;	14'h2938: data <= 32'hC89C89C9;	14'h2939: data <= 32'hC84B48CC;	14'h293A: data <= 32'hC7FA07CF;	14'h293B: data <= 32'hC7A8C6D2;	14'h293C: data <= 32'hC75785D5;	14'h293D: data <= 32'hC6FBD49D;	14'h293E: data <= 32'hC67FA9C7;	14'h293F: data <= 32'hC6037EF1;	14'h2940: data <= 32'hC587541B;	14'h2941: data <= 32'hC50B2945;	14'h2942: data <= 32'hC48EFE6F;	14'h2943: data <= 32'hC412D399;	14'h2944: data <= 32'hC396A8C3;	14'h2945: data <= 32'hC31A7DED;	14'h2946: data <= 32'hC29E5317;	14'h2947: data <= 32'hC2222841;	14'h2948: data <= 32'hC1A5FD6B;	14'h2949: data <= 32'hC129D295;	14'h294A: data <= 32'hC0ADA7BF;	14'h294B: data <= 32'hC0317CE9;	14'h294C: data <= 32'hBFB55213;	14'h294D: data <= 32'hBF38EFC5;	14'h294E: data <= 32'hBEB4C0A1;	14'h294F: data <= 32'hBE30917D;	14'h2950: data <= 32'hBDAC6259;	14'h2951: data <= 32'hBD283335;	14'h2952: data <= 32'hBCA40410;	14'h2953: data <= 32'hBC1FD4EC;	14'h2954: data <= 32'hBB9BA5C8;	14'h2955: data <= 32'hBB1776A4;	14'h2956: data <= 32'hBA934780;	14'h2957: data <= 32'hBA0F185B;	14'h2958: data <= 32'hB98AE937;	14'h2959: data <= 32'hB906BA13;	14'h295A: data <= 32'hB8828AEF;	14'h295B: data <= 32'hB7FE5BCB;	14'h295C: data <= 32'hB77A2CA7;	14'h295D: data <= 32'hB6F5FD82;	14'h295E: data <= 32'hB6492DB0;	14'h295F: data <= 32'hB592E309;	14'h2960: data <= 32'hB4DC9863;	14'h2961: data <= 32'hB4264DBD;	14'h2962: data <= 32'hB3700317;	14'h2963: data <= 32'hB2B9B871;	14'h2964: data <= 32'hB2036DCB;	14'h2965: data <= 32'hB14D2324;	14'h2966: data <= 32'hB096D87E;	14'h2967: data <= 32'hAFE08DD8;	14'h2968: data <= 32'hAF2A4332;	14'h2969: data <= 32'hAE73F88C;	14'h296A: data <= 32'hADBDADE5;	14'h296B: data <= 32'hAD07633F;	14'h296C: data <= 32'hAC511899;	14'h296D: data <= 32'hAB9ACDF3;	14'h296E: data <= 32'hA9BA4F35;	14'h296F: data <= 32'hA70E7E66;	14'h2970: data <= 32'hA462AD98;	14'h2971: data <= 32'hA1B6DCC9;	14'h2972: data <= 32'h9F0B0BFB;	14'h2973: data <= 32'h9C5F3B2C;	14'h2974: data <= 32'h99B36A5E;	14'h2975: data <= 32'h9707998F;	14'h2976: data <= 32'h945BC8C1;	14'h2977: data <= 32'h91AFF7F2;	14'h2978: data <= 32'h8F042724;	14'h2979: data <= 32'h8C585655;	14'h297A: data <= 32'h89AC8587;	14'h297B: data <= 32'h8700B4B8;	14'h297C: data <= 32'h8454E3EA;	14'h297D: data <= 32'h81A9131B;	14'h297E: data <= 32'h80E06587;	14'h297F: data <= 32'h833171D3;	14'h2980: data <= 32'h85827E1F;	14'h2981: data <= 32'h87D38A6A;	14'h2982: data <= 32'h8A2496B6;	14'h2983: data <= 32'h8C75A302;	14'h2984: data <= 32'h8EC6AF4E;	14'h2985: data <= 32'h9117BB9A;	14'h2986: data <= 32'h9368C7E6;	14'h2987: data <= 32'h95B9D432;	14'h2988: data <= 32'h980AE07D;	14'h2989: data <= 32'h9A5BECC9;	14'h298A: data <= 32'h9CACF915;	14'h298B: data <= 32'h9EFE0561;	14'h298C: data <= 32'hA14F11AD;	14'h298D: data <= 32'hA3A01DF9;	14'h298E: data <= 32'hA5B41F8D;	14'h298F: data <= 32'hA68CBF1A;	14'h2990: data <= 32'hA7655EA7;	14'h2991: data <= 32'hA83DFE35;	14'h2992: data <= 32'hA9169DC2;	14'h2993: data <= 32'hA9EF3D4F;	14'h2994: data <= 32'hAAC7DCDC;	14'h2995: data <= 32'hABA07C69;	14'h2996: data <= 32'hAC791BF6;	14'h2997: data <= 32'hAD51BB83;	14'h2998: data <= 32'hAE2A5B10;	14'h2999: data <= 32'hAF02FA9D;	14'h299A: data <= 32'hAFDB9A2A;	14'h299B: data <= 32'hB0B439B7;	14'h299C: data <= 32'hB18CD944;	14'h299D: data <= 32'hB26578D1;	14'h299E: data <= 32'hB33E185F;	14'h299F: data <= 32'hB3DAB088;	14'h29A0: data <= 32'hB473DA8F;	14'h29A1: data <= 32'hB50D0496;	14'h29A2: data <= 32'hB5A62E9D;	14'h29A3: data <= 32'hB63F58A4;	14'h29A4: data <= 32'hB6D882AA;	14'h29A5: data <= 32'hB771ACB1;	14'h29A6: data <= 32'hB80AD6B8;	14'h29A7: data <= 32'hB8A400BF;	14'h29A8: data <= 32'hB93D2AC6;	14'h29A9: data <= 32'hB9D654CC;	14'h29AA: data <= 32'hBA6F7ED3;	14'h29AB: data <= 32'hBB08A8DA;	14'h29AC: data <= 32'hBBA1D2E1;	14'h29AD: data <= 32'hBC3AFCE8;	14'h29AE: data <= 32'hBCD426EF;	14'h29AF: data <= 32'hBD64BF83;	14'h29B0: data <= 32'hBDF22BB4;	14'h29B1: data <= 32'hBE7F97E4;	14'h29B2: data <= 32'hBF0D0415;	14'h29B3: data <= 32'hBF9A7046;	14'h29B4: data <= 32'hC027DC77;	14'h29B5: data <= 32'hC0B548A8;	14'h29B6: data <= 32'hC142B4D8;	14'h29B7: data <= 32'hC1D02109;	14'h29B8: data <= 32'hC25D8D3A;	14'h29B9: data <= 32'hC2EAF96B;	14'h29BA: data <= 32'hC378659C;	14'h29BB: data <= 32'hC405D1CD;	14'h29BC: data <= 32'hC4933DFD;	14'h29BD: data <= 32'hC520AA2E;	14'h29BE: data <= 32'hC5AE165F;	14'h29BF: data <= 32'hC61F815B;	14'h29C0: data <= 32'hC6766475;	14'h29C1: data <= 32'hC6CD478F;	14'h29C2: data <= 32'hC7242AA9;	14'h29C3: data <= 32'hC77B0DC3;	14'h29C4: data <= 32'hC7D1F0DD;	14'h29C5: data <= 32'hC828D3F8;	14'h29C6: data <= 32'hC87FB712;	14'h29C7: data <= 32'hC8D69A2C;	14'h29C8: data <= 32'hC92D7D46;	14'h29C9: data <= 32'hC9846060;	14'h29CA: data <= 32'hC9DB437A;	14'h29CB: data <= 32'hCA322694;	14'h29CC: data <= 32'hCA8909AE;	14'h29CD: data <= 32'hCADFECC9;	14'h29CE: data <= 32'hCB36CFE3;	14'h29CF: data <= 32'hCB7CC22F;	14'h29D0: data <= 32'hCB9AA9D9;	14'h29D1: data <= 32'hCBB89183;	14'h29D2: data <= 32'hCBD6792D;	14'h29D3: data <= 32'hCBF460D8;	14'h29D4: data <= 32'hCC124882;	14'h29D5: data <= 32'hCC30302C;	14'h29D6: data <= 32'hCC4E17D6;	14'h29D7: data <= 32'hCC6BFF80;	14'h29D8: data <= 32'hCC89E72B;	14'h29D9: data <= 32'hCCA7CED5;	14'h29DA: data <= 32'hCCC5B67F;	14'h29DB: data <= 32'hCCE39E29;	14'h29DC: data <= 32'hCD0185D4;	14'h29DD: data <= 32'hCD1F6D7E;	14'h29DE: data <= 32'hCD3D5528;	14'h29DF: data <= 32'hCD59AD2D;	14'h29E0: data <= 32'hCD6453DF;	14'h29E1: data <= 32'hCD6EFA91;	14'h29E2: data <= 32'hCD79A143;	14'h29E3: data <= 32'hCD8447F5;	14'h29E4: data <= 32'hCD8EEEA7;	14'h29E5: data <= 32'hCD999559;	14'h29E6: data <= 32'hCDA43C0B;	14'h29E7: data <= 32'hCDAEE2BD;	14'h29E8: data <= 32'hCDB9896F;	14'h29E9: data <= 32'hCDC43021;	14'h29EA: data <= 32'hCDCED6D3;	14'h29EB: data <= 32'hCDD97D85;	14'h29EC: data <= 32'hCDE42437;	14'h29ED: data <= 32'hCDEECAE9;	14'h29EE: data <= 32'hCDF9719B;	14'h29EF: data <= 32'hCE04184D;	14'h29F0: data <= 32'hCE12C38E;	14'h29F1: data <= 32'hCE220F85;	14'h29F2: data <= 32'hCE315B7C;	14'h29F3: data <= 32'hCE40A774;	14'h29F4: data <= 32'hCE4FF36B;	14'h29F5: data <= 32'hCE5F3F62;	14'h29F6: data <= 32'hCE6E8B5A;	14'h29F7: data <= 32'hCE7DD751;	14'h29F8: data <= 32'hCE8D2349;	14'h29F9: data <= 32'hCE9C6F40;	14'h29FA: data <= 32'hCEABBB37;	14'h29FB: data <= 32'hCEBB072F;	14'h29FC: data <= 32'hCECA5326;	14'h29FD: data <= 32'hCED99F1D;	14'h29FE: data <= 32'hCEE8EB15;	14'h29FF: data <= 32'hCEF8370C;	14'h2A00: data <= 32'hCF086AFA;	14'h2A01: data <= 32'hCF191C8C;	14'h2A02: data <= 32'hCF29CE1F;	14'h2A03: data <= 32'hCF3A7FB2;	14'h2A04: data <= 32'hCF4B3144;	14'h2A05: data <= 32'hCF5BE2D7;	14'h2A06: data <= 32'hCF6C946A;	14'h2A07: data <= 32'hCF7D45FC;	14'h2A08: data <= 32'hCF8DF78F;	14'h2A09: data <= 32'hCF9EA922;	14'h2A0A: data <= 32'hCFAF5AB4;	14'h2A0B: data <= 32'hCFC00C47;	14'h2A0C: data <= 32'hCFD0BDDA;	14'h2A0D: data <= 32'hCFE16F6D;	14'h2A0E: data <= 32'hCFF220FF;	14'h2A0F: data <= 32'hD002D292;	14'h2A10: data <= 32'hD01A3A66;	14'h2A11: data <= 32'hD03A716E;	14'h2A12: data <= 32'hD05AA877;	14'h2A13: data <= 32'hD07ADF80;	14'h2A14: data <= 32'hD09B1689;	14'h2A15: data <= 32'hD0BB4D92;	14'h2A16: data <= 32'hD0DB849B;	14'h2A17: data <= 32'hD0FBBBA4;	14'h2A18: data <= 32'hD11BF2AD;	14'h2A19: data <= 32'hD13C29B6;	14'h2A1A: data <= 32'hD15C60BF;	14'h2A1B: data <= 32'hD17C97C7;	14'h2A1C: data <= 32'hD19CCED0;	14'h2A1D: data <= 32'hD1BD05D9;	14'h2A1E: data <= 32'hD1DD3CE2;	14'h2A1F: data <= 32'hD1FD73EB;	14'h2A20: data <= 32'hD22092ED;	14'h2A21: data <= 32'hD24E3AD7;	14'h2A22: data <= 32'hD27BE2C0;	14'h2A23: data <= 32'hD2A98AA9;	14'h2A24: data <= 32'hD2D73293;	14'h2A25: data <= 32'hD304DA7C;	14'h2A26: data <= 32'hD3328266;	14'h2A27: data <= 32'hD3602A4F;	14'h2A28: data <= 32'hD38DD238;	14'h2A29: data <= 32'hD3BB7A22;	14'h2A2A: data <= 32'hD3E9220B;	14'h2A2B: data <= 32'hD416C9F5;	14'h2A2C: data <= 32'hD44471DE;	14'h2A2D: data <= 32'hD47219C7;	14'h2A2E: data <= 32'hD49FC1B1;	14'h2A2F: data <= 32'hD4CD699A;	14'h2A30: data <= 32'hD4FB1183;	14'h2A31: data <= 32'hD51FDD7E;	14'h2A32: data <= 32'hD544A978;	14'h2A33: data <= 32'hD5697572;	14'h2A34: data <= 32'hD58E416C;	14'h2A35: data <= 32'hD5B30D66;	14'h2A36: data <= 32'hD5D7D960;	14'h2A37: data <= 32'hD5FCA55A;	14'h2A38: data <= 32'hD6217154;	14'h2A39: data <= 32'hD6463D4E;	14'h2A3A: data <= 32'hD66B0948;	14'h2A3B: data <= 32'hD68FD543;	14'h2A3C: data <= 32'hD6B4A13D;	14'h2A3D: data <= 32'hD6D96D37;	14'h2A3E: data <= 32'hD6FE3931;	14'h2A3F: data <= 32'hD723052B;	14'h2A40: data <= 32'hD747D125;	14'h2A41: data <= 32'hD75F09F0;	14'h2A42: data <= 32'hD772840F;	14'h2A43: data <= 32'hD785FE2E;	14'h2A44: data <= 32'hD799784D;	14'h2A45: data <= 32'hD7ACF26C;	14'h2A46: data <= 32'hD7C06C8B;	14'h2A47: data <= 32'hD7D3E6AB;	14'h2A48: data <= 32'hD7E760CA;	14'h2A49: data <= 32'hD7FADAE9;	14'h2A4A: data <= 32'hD80E5508;	14'h2A4B: data <= 32'hD821CF27;	14'h2A4C: data <= 32'hD8354946;	14'h2A4D: data <= 32'hD848C365;	14'h2A4E: data <= 32'hD85C3D84;	14'h2A4F: data <= 32'hD86FB7A3;	14'h2A50: data <= 32'hD88331C2;	14'h2A51: data <= 32'hD8919C0A;	14'h2A52: data <= 32'hD89C2B04;	14'h2A53: data <= 32'hD8A6B9FE;	14'h2A54: data <= 32'hD8B148F7;	14'h2A55: data <= 32'hD8BBD7F1;	14'h2A56: data <= 32'hD8C666EA;	14'h2A57: data <= 32'hD8D0F5E4;	14'h2A58: data <= 32'hD8DB84DE;	14'h2A59: data <= 32'hD8E613D7;	14'h2A5A: data <= 32'hD8F0A2D1;	14'h2A5B: data <= 32'hD8FB31CB;	14'h2A5C: data <= 32'hD905C0C4;	14'h2A5D: data <= 32'hD9104FBE;	14'h2A5E: data <= 32'hD91ADEB7;	14'h2A5F: data <= 32'hD9256DB1;	14'h2A60: data <= 32'hD92FFCAB;	14'h2A61: data <= 32'hD93A3441;	14'h2A62: data <= 32'hD943CA83;	14'h2A63: data <= 32'hD94D60C5;	14'h2A64: data <= 32'hD956F707;	14'h2A65: data <= 32'hD9608D49;	14'h2A66: data <= 32'hD96A238B;	14'h2A67: data <= 32'hD973B9CD;	14'h2A68: data <= 32'hD97D500F;	14'h2A69: data <= 32'hD986E651;	14'h2A6A: data <= 32'hD9907C93;	14'h2A6B: data <= 32'hD99A12D5;	14'h2A6C: data <= 32'hD9A3A917;	14'h2A6D: data <= 32'hD9AD3F59;	14'h2A6E: data <= 32'hD9B6D59B;	14'h2A6F: data <= 32'hD9C06BDD;	14'h2A70: data <= 32'hD9CA0220;	14'h2A71: data <= 32'hD9D37479;	14'h2A72: data <= 32'hD9DC00FF;	14'h2A73: data <= 32'hD9E48D85;	14'h2A74: data <= 32'hD9ED1A0B;	14'h2A75: data <= 32'hD9F5A691;	14'h2A76: data <= 32'hD9FE3317;	14'h2A77: data <= 32'hDA06BF9D;	14'h2A78: data <= 32'hDA0F4C23;	14'h2A79: data <= 32'hDA17D8A9;	14'h2A7A: data <= 32'hDA20652F;	14'h2A7B: data <= 32'hDA28F1B5;	14'h2A7C: data <= 32'hDA317E3B;	14'h2A7D: data <= 32'hDA3A0AC2;	14'h2A7E: data <= 32'hDA429748;	14'h2A7F: data <= 32'hDA4B23CE;	14'h2A80: data <= 32'hDA53B054;	14'h2A81: data <= 32'hDA5C3CDA;	14'h2A82: data <= 32'hDA6E0C93;	14'h2A83: data <= 32'hDA80AD84;	14'h2A84: data <= 32'hDA934E76;	14'h2A85: data <= 32'hDAA5EF68;	14'h2A86: data <= 32'hDAB8905A;	14'h2A87: data <= 32'hDACB314C;	14'h2A88: data <= 32'hDADDD23E;	14'h2A89: data <= 32'hDAF07330;	14'h2A8A: data <= 32'hDB031422;	14'h2A8B: data <= 32'hDB15B514;	14'h2A8C: data <= 32'hDB285606;	14'h2A8D: data <= 32'hDB3AF6F8;	14'h2A8E: data <= 32'hDB4D97E9;	14'h2A8F: data <= 32'hDB6038DB;	14'h2A90: data <= 32'hDB72D9CD;	14'h2A91: data <= 32'hDB857ABF;	14'h2A92: data <= 32'hDB9C7AA2;	14'h2A93: data <= 32'hDBB553EC;	14'h2A94: data <= 32'hDBCE2D35;	14'h2A95: data <= 32'hDBE7067E;	14'h2A96: data <= 32'hDBFFDFC7;	14'h2A97: data <= 32'hDC18B911;	14'h2A98: data <= 32'hDC31925A;	14'h2A99: data <= 32'hDC4A6BA3;	14'h2A9A: data <= 32'hDC6344EC;	14'h2A9B: data <= 32'hDC7C1E36;	14'h2A9C: data <= 32'hDC94F77F;	14'h2A9D: data <= 32'hDCADD0C8;	14'h2A9E: data <= 32'hDCC6AA11;	14'h2A9F: data <= 32'hDCDF835B;	14'h2AA0: data <= 32'hDCF85CA4;	14'h2AA1: data <= 32'hDD1135ED;	14'h2AA2: data <= 32'hDD28A0B5;	14'h2AA3: data <= 32'hDD3E889F;	14'h2AA4: data <= 32'hDD54708A;	14'h2AA5: data <= 32'hDD6A5874;	14'h2AA6: data <= 32'hDD80405E;	14'h2AA7: data <= 32'hDD962848;	14'h2AA8: data <= 32'hDDAC1033;	14'h2AA9: data <= 32'hDDC1F81D;	14'h2AAA: data <= 32'hDDD7E007;	14'h2AAB: data <= 32'hDDEDC7F1;	14'h2AAC: data <= 32'hDE03AFDB;	14'h2AAD: data <= 32'hDE1997C6;	14'h2AAE: data <= 32'hDE2F7FB0;	14'h2AAF: data <= 32'hDE45679A;	14'h2AB0: data <= 32'hDE5B4F84;	14'h2AB1: data <= 32'hDE71376E;	14'h2AB2: data <= 32'hDE86D87A;	14'h2AB3: data <= 32'hDE9BBA2F;	14'h2AB4: data <= 32'hDEB09BE3;	14'h2AB5: data <= 32'hDEC57D98;	14'h2AB6: data <= 32'hDEDA5F4C;	14'h2AB7: data <= 32'hDEEF4100;	14'h2AB8: data <= 32'hDF0422B5;	14'h2AB9: data <= 32'hDF190469;	14'h2ABA: data <= 32'hDF2DE61D;	14'h2ABB: data <= 32'hDF42C7D2;	14'h2ABC: data <= 32'hDF57A986;	14'h2ABD: data <= 32'hDF6C8B3B;	14'h2ABE: data <= 32'hDF816CEF;	14'h2ABF: data <= 32'hDF964EA3;	14'h2AC0: data <= 32'hDFAB3058;	14'h2AC1: data <= 32'hDFC0120C;	14'h2AC2: data <= 32'hDFD4B629;	14'h2AC3: data <= 32'hDFE52471;	14'h2AC4: data <= 32'hDFF592B9;	14'h2AC5: data <= 32'hE0060100;	14'h2AC6: data <= 32'hE0166F48;	14'h2AC7: data <= 32'hE026DD90;	14'h2AC8: data <= 32'hE0374BD7;	14'h2AC9: data <= 32'hE047BA1F;	14'h2ACA: data <= 32'hE0582867;	14'h2ACB: data <= 32'hE06896AE;	14'h2ACC: data <= 32'hE07904F6;	14'h2ACD: data <= 32'hE089733E;	14'h2ACE: data <= 32'hE099E185;	14'h2ACF: data <= 32'hE0AA4FCD;	14'h2AD0: data <= 32'hE0BABE15;	14'h2AD1: data <= 32'hE0CB2C5C;	14'h2AD2: data <= 32'hE0DB9AA4;	14'h2AD3: data <= 32'hE0E9266E;	14'h2AD4: data <= 32'hE0F62349;	14'h2AD5: data <= 32'hE1032023;	14'h2AD6: data <= 32'hE1101CFE;	14'h2AD7: data <= 32'hE11D19D9;	14'h2AD8: data <= 32'hE12A16B4;	14'h2AD9: data <= 32'hE137138E;	14'h2ADA: data <= 32'hE1441069;	14'h2ADB: data <= 32'hE1510D44;	14'h2ADC: data <= 32'hE15E0A1E;	14'h2ADD: data <= 32'hE16B06F9;	14'h2ADE: data <= 32'hE17803D4;	14'h2ADF: data <= 32'hE18500AF;	14'h2AE0: data <= 32'hE191FD89;	14'h2AE1: data <= 32'hE19EFA64;	14'h2AE2: data <= 32'hE1ABF73F;	14'h2AE3: data <= 32'hE1B7FB41;	14'h2AE4: data <= 32'hE1C367CA;	14'h2AE5: data <= 32'hE1CED452;	14'h2AE6: data <= 32'hE1DA40DB;	14'h2AE7: data <= 32'hE1E5AD64;	14'h2AE8: data <= 32'hE1F119ED;	14'h2AE9: data <= 32'hE1FC8676;	14'h2AEA: data <= 32'hE207F2FF;	14'h2AEB: data <= 32'hE2135F88;	14'h2AEC: data <= 32'hE21ECC11;	14'h2AED: data <= 32'hE22A389A;	14'h2AEE: data <= 32'hE235A522;	14'h2AEF: data <= 32'hE24111AB;	14'h2AF0: data <= 32'hE24C7E34;	14'h2AF1: data <= 32'hE257EABD;	14'h2AF2: data <= 32'hE2635746;	14'h2AF3: data <= 32'hE26E94FB;	14'h2AF4: data <= 32'hE2798E02;	14'h2AF5: data <= 32'hE284870A;	14'h2AF6: data <= 32'hE28F8011;	14'h2AF7: data <= 32'hE29A7918;	14'h2AF8: data <= 32'hE2A5721F;	14'h2AF9: data <= 32'hE2B06B26;	14'h2AFA: data <= 32'hE2BB642E;	14'h2AFB: data <= 32'hE2C65D35;	14'h2AFC: data <= 32'hE2D1563C;	14'h2AFD: data <= 32'hE2DC4F43;	14'h2AFE: data <= 32'hE2E7484A;	14'h2AFF: data <= 32'hE2F24152;	14'h2B00: data <= 32'hE2FD3A59;	14'h2B01: data <= 32'hE3083360;	14'h2B02: data <= 32'hE3132C67;	14'h2B03: data <= 32'hE31EA379;	14'h2B04: data <= 32'hE32C36BA;	14'h2B05: data <= 32'hE339C9FB;	14'h2B06: data <= 32'hE3475D3C;	14'h2B07: data <= 32'hE354F07D;	14'h2B08: data <= 32'hE36283BE;	14'h2B09: data <= 32'hE37016FF;	14'h2B0A: data <= 32'hE37DAA40;	14'h2B0B: data <= 32'hE38B3D81;	14'h2B0C: data <= 32'hE398D0C2;	14'h2B0D: data <= 32'hE3A66403;	14'h2B0E: data <= 32'hE3B3F744;	14'h2B0F: data <= 32'hE3C18A85;	14'h2B10: data <= 32'hE3CF1DC6;	14'h2B11: data <= 32'hE3DCB107;	14'h2B12: data <= 32'hE3EA4448;	14'h2B13: data <= 32'hE3F7D789;	14'h2B14: data <= 32'hE406353B;	14'h2B15: data <= 32'hE414988D;	14'h2B16: data <= 32'hE422FBDF;	14'h2B17: data <= 32'hE4315F31;	14'h2B18: data <= 32'hE43FC283;	14'h2B19: data <= 32'hE44E25D5;	14'h2B1A: data <= 32'hE45C8927;	14'h2B1B: data <= 32'hE46AEC79;	14'h2B1C: data <= 32'hE4794FCB;	14'h2B1D: data <= 32'hE487B31D;	14'h2B1E: data <= 32'hE496166F;	14'h2B1F: data <= 32'hE4A479C1;	14'h2B20: data <= 32'hE4B2DD13;	14'h2B21: data <= 32'hE4C14065;	14'h2B22: data <= 32'hE4CFA3B7;	14'h2B23: data <= 32'hE4DE0709;	14'h2B24: data <= 32'hE4E95573;	14'h2B25: data <= 32'hE4F3A64A;	14'h2B26: data <= 32'hE4FDF721;	14'h2B27: data <= 32'hE50847F8;	14'h2B28: data <= 32'hE51298CE;	14'h2B29: data <= 32'hE51CE9A5;	14'h2B2A: data <= 32'hE5273A7C;	14'h2B2B: data <= 32'hE5318B52;	14'h2B2C: data <= 32'hE53BDC29;	14'h2B2D: data <= 32'hE5462D00;	14'h2B2E: data <= 32'hE5507DD6;	14'h2B2F: data <= 32'hE55ACEAD;	14'h2B30: data <= 32'hE5651F84;	14'h2B31: data <= 32'hE56F705A;	14'h2B32: data <= 32'hE579C131;	14'h2B33: data <= 32'hE5841208;	14'h2B34: data <= 32'hE58CAAD8;	14'h2B35: data <= 32'hE593CDA3;	14'h2B36: data <= 32'hE59AF06E;	14'h2B37: data <= 32'hE5A21338;	14'h2B38: data <= 32'hE5A93603;	14'h2B39: data <= 32'hE5B058CE;	14'h2B3A: data <= 32'hE5B77B99;	14'h2B3B: data <= 32'hE5BE9E64;	14'h2B3C: data <= 32'hE5C5C12E;	14'h2B3D: data <= 32'hE5CCE3F9;	14'h2B3E: data <= 32'hE5D406C4;	14'h2B3F: data <= 32'hE5DB298F;	14'h2B40: data <= 32'hE5E24C59;	14'h2B41: data <= 32'hE5E96F24;	14'h2B42: data <= 32'hE5F091EF;	14'h2B43: data <= 32'hE5F7B4BA;	14'h2B44: data <= 32'hE5FEFD09;	14'h2B45: data <= 32'hE6069382;	14'h2B46: data <= 32'hE60E29FA;	14'h2B47: data <= 32'hE615C072;	14'h2B48: data <= 32'hE61D56EB;	14'h2B49: data <= 32'hE624ED63;	14'h2B4A: data <= 32'hE62C83DC;	14'h2B4B: data <= 32'hE6341A54;	14'h2B4C: data <= 32'hE63BB0CD;	14'h2B4D: data <= 32'hE6434745;	14'h2B4E: data <= 32'hE64ADDBE;	14'h2B4F: data <= 32'hE6527436;	14'h2B50: data <= 32'hE65A0AAF;	14'h2B51: data <= 32'hE661A127;	14'h2B52: data <= 32'hE66937A0;	14'h2B53: data <= 32'hE670CE18;	14'h2B54: data <= 32'hE678E8DF;	14'h2B55: data <= 32'hE6854729;	14'h2B56: data <= 32'hE691A574;	14'h2B57: data <= 32'hE69E03BE;	14'h2B58: data <= 32'hE6AA6208;	14'h2B59: data <= 32'hE6B6C053;	14'h2B5A: data <= 32'hE6C31E9D;	14'h2B5B: data <= 32'hE6CF7CE8;	14'h2B5C: data <= 32'hE6DBDB32;	14'h2B5D: data <= 32'hE6E8397C;	14'h2B5E: data <= 32'hE6F497C7;	14'h2B5F: data <= 32'hE700F611;	14'h2B60: data <= 32'hE70D545C;	14'h2B61: data <= 32'hE719B2A6;	14'h2B62: data <= 32'hE72610F0;	14'h2B63: data <= 32'hE7326F3B;	14'h2B64: data <= 32'hE73ECD85;	14'h2B65: data <= 32'hE74C825E;	14'h2B66: data <= 32'hE75A60BC;	14'h2B67: data <= 32'hE7683F1A;	14'h2B68: data <= 32'hE7761D78;	14'h2B69: data <= 32'hE783FBD6;	14'h2B6A: data <= 32'hE791DA34;	14'h2B6B: data <= 32'hE79FB892;	14'h2B6C: data <= 32'hE7AD96F0;	14'h2B6D: data <= 32'hE7BB754E;	14'h2B6E: data <= 32'hE7C953AD;	14'h2B6F: data <= 32'hE7D7320B;	14'h2B70: data <= 32'hE7E51069;	14'h2B71: data <= 32'hE7F2EEC7;	14'h2B72: data <= 32'hE800CD25;	14'h2B73: data <= 32'hE80EAB83;	14'h2B74: data <= 32'hE81C89E1;	14'h2B75: data <= 32'hE8275290;	14'h2B76: data <= 32'hE830A033;	14'h2B77: data <= 32'hE839EDD6;	14'h2B78: data <= 32'hE8433B79;	14'h2B79: data <= 32'hE84C891C;	14'h2B7A: data <= 32'hE855D6BF;	14'h2B7B: data <= 32'hE85F2462;	14'h2B7C: data <= 32'hE8687204;	14'h2B7D: data <= 32'hE871BFA7;	14'h2B7E: data <= 32'hE87B0D4A;	14'h2B7F: data <= 32'hE8845AED;	14'h2B80: data <= 32'hE88DA890;	14'h2B81: data <= 32'hE896F633;	14'h2B82: data <= 32'hE8A043D6;	14'h2B83: data <= 32'hE8A99179;	14'h2B84: data <= 32'hE8B2DF1C;	14'h2B85: data <= 32'hE8B9CEE5;	14'h2B86: data <= 32'hE8BDF5EA;	14'h2B87: data <= 32'hE8C21CF0;	14'h2B88: data <= 32'hE8C643F6;	14'h2B89: data <= 32'hE8CA6AFB;	14'h2B8A: data <= 32'hE8CE9201;	14'h2B8B: data <= 32'hE8D2B906;	14'h2B8C: data <= 32'hE8D6E00C;	14'h2B8D: data <= 32'hE8DB0712;	14'h2B8E: data <= 32'hE8DF2E17;	14'h2B8F: data <= 32'hE8E3551D;	14'h2B90: data <= 32'hE8E77C22;	14'h2B91: data <= 32'hE8EBA328;	14'h2B92: data <= 32'hE8EFCA2D;	14'h2B93: data <= 32'hE8F3F133;	14'h2B94: data <= 32'hE8F81839;	14'h2B95: data <= 32'hE8FC2159;	14'h2B96: data <= 32'hE8FFCD79;	14'h2B97: data <= 32'hE9037999;	14'h2B98: data <= 32'hE90725B9;	14'h2B99: data <= 32'hE90AD1D9;	14'h2B9A: data <= 32'hE90E7DF8;	14'h2B9B: data <= 32'hE9122A18;	14'h2B9C: data <= 32'hE915D638;	14'h2B9D: data <= 32'hE9198258;	14'h2B9E: data <= 32'hE91D2E78;	14'h2B9F: data <= 32'hE920DA97;	14'h2BA0: data <= 32'hE92486B7;	14'h2BA1: data <= 32'hE92832D7;	14'h2BA2: data <= 32'hE92BDEF7;	14'h2BA3: data <= 32'hE92F8B17;	14'h2BA4: data <= 32'hE9333736;	14'h2BA5: data <= 32'hE936E810;	14'h2BA6: data <= 32'hE93B42FE;	14'h2BA7: data <= 32'hE93F9DEC;	14'h2BA8: data <= 32'hE943F8DB;	14'h2BA9: data <= 32'hE94853C9;	14'h2BAA: data <= 32'hE94CAEB7;	14'h2BAB: data <= 32'hE95109A6;	14'h2BAC: data <= 32'hE9556494;	14'h2BAD: data <= 32'hE959BF82;	14'h2BAE: data <= 32'hE95E1A70;	14'h2BAF: data <= 32'hE962755F;	14'h2BB0: data <= 32'hE966D04D;	14'h2BB1: data <= 32'hE96B2B3B;	14'h2BB2: data <= 32'hE96F862A;	14'h2BB3: data <= 32'hE973E118;	14'h2BB4: data <= 32'hE9783C06;	14'h2BB5: data <= 32'hE97C96F5;	14'h2BB6: data <= 32'hE98025B7;	14'h2BB7: data <= 32'hE98384D6;	14'h2BB8: data <= 32'hE986E3F5;	14'h2BB9: data <= 32'hE98A4313;	14'h2BBA: data <= 32'hE98DA232;	14'h2BBB: data <= 32'hE9910151;	14'h2BBC: data <= 32'hE994606F;	14'h2BBD: data <= 32'hE997BF8E;	14'h2BBE: data <= 32'hE99B1EAD;	14'h2BBF: data <= 32'hE99E7DCB;	14'h2BC0: data <= 32'hE9A1DCEA;	14'h2BC1: data <= 32'hE9A53C09;	14'h2BC2: data <= 32'hE9A89B28;	14'h2BC3: data <= 32'hE9ABFA46;	14'h2BC4: data <= 32'hE9AF5965;	14'h2BC5: data <= 32'hE9B2B884;	14'h2BC6: data <= 32'hE9B6296B;	14'h2BC7: data <= 32'hE9B9A672;	14'h2BC8: data <= 32'hE9BD2379;	14'h2BC9: data <= 32'hE9C0A080;	14'h2BCA: data <= 32'hE9C41D87;	14'h2BCB: data <= 32'hE9C79A8E;	14'h2BCC: data <= 32'hE9CB1795;	14'h2BCD: data <= 32'hE9CE949D;	14'h2BCE: data <= 32'hE9D211A4;	14'h2BCF: data <= 32'hE9D58EAB;	14'h2BD0: data <= 32'hE9D90BB2;	14'h2BD1: data <= 32'hE9DC88B9;	14'h2BD2: data <= 32'hE9E005C0;	14'h2BD3: data <= 32'hE9E382C7;	14'h2BD4: data <= 32'hE9E6FFCE;	14'h2BD5: data <= 32'hE9EA7CD5;	14'h2BD6: data <= 32'hE9ECDAF3;	14'h2BD7: data <= 32'hE9ED61B5;	14'h2BD8: data <= 32'hE9EDE877;	14'h2BD9: data <= 32'hE9EE6F39;	14'h2BDA: data <= 32'hE9EEF5FB;	14'h2BDB: data <= 32'hE9EF7CBC;	14'h2BDC: data <= 32'hE9F0037E;	14'h2BDD: data <= 32'hE9F08A40;	14'h2BDE: data <= 32'hE9F11102;	14'h2BDF: data <= 32'hE9F197C4;	14'h2BE0: data <= 32'hE9F21E86;	14'h2BE1: data <= 32'hE9F2A548;	14'h2BE2: data <= 32'hE9F32C0A;	14'h2BE3: data <= 32'hE9F3B2CC;	14'h2BE4: data <= 32'hE9F4398E;	14'h2BE5: data <= 32'hE9F4C050;	14'h2BE6: data <= 32'hE9F540DE;	14'h2BE7: data <= 32'hE9F5A162;	14'h2BE8: data <= 32'hE9F601E5;	14'h2BE9: data <= 32'hE9F66268;	14'h2BEA: data <= 32'hE9F6C2EC;	14'h2BEB: data <= 32'hE9F7236F;	14'h2BEC: data <= 32'hE9F783F3;	14'h2BED: data <= 32'hE9F7E476;	14'h2BEE: data <= 32'hE9F844FA;	14'h2BEF: data <= 32'hE9F8A57D;	14'h2BF0: data <= 32'hE9F90600;	14'h2BF1: data <= 32'hE9F96684;	14'h2BF2: data <= 32'hE9F9C707;	14'h2BF3: data <= 32'hE9FA278B;	14'h2BF4: data <= 32'hE9FA880E;	14'h2BF5: data <= 32'hE9FAE892;	14'h2BF6: data <= 32'hE9FB4915;	14'h2BF7: data <= 32'hE9FEB58F;	14'h2BF8: data <= 32'hEA024E9A;	14'h2BF9: data <= 32'hEA05E7A6;	14'h2BFA: data <= 32'hEA0980B1;	14'h2BFB: data <= 32'hEA0D19BD;	14'h2BFC: data <= 32'hEA10B2C8;	14'h2BFD: data <= 32'hEA144BD4;	14'h2BFE: data <= 32'hEA17E4DF;	14'h2BFF: data <= 32'hEA1B7DEB;	14'h2C00: data <= 32'hEA1F16F6;	14'h2C01: data <= 32'hEA22B002;	14'h2C02: data <= 32'hEA26490D;	14'h2C03: data <= 32'hEA29E219;	14'h2C04: data <= 32'hEA2D7B24;	14'h2C05: data <= 32'hEA311430;	14'h2C06: data <= 32'hEA34AD3B;	14'h2C07: data <= 32'hEA36626F;	14'h2C08: data <= 32'hEA37646E;	14'h2C09: data <= 32'hEA38666E;	14'h2C0A: data <= 32'hEA39686E;	14'h2C0B: data <= 32'hEA3A6A6E;	14'h2C0C: data <= 32'hEA3B6C6D;	14'h2C0D: data <= 32'hEA3C6E6D;	14'h2C0E: data <= 32'hEA3D706D;	14'h2C0F: data <= 32'hEA3E726D;	14'h2C10: data <= 32'hEA3F746C;	14'h2C11: data <= 32'hEA40766C;	14'h2C12: data <= 32'hEA41786C;	14'h2C13: data <= 32'hEA427A6C;	14'h2C14: data <= 32'hEA437C6C;	14'h2C15: data <= 32'hEA447E6B;	14'h2C16: data <= 32'hEA45806B;	14'h2C17: data <= 32'hEA453570;	14'h2C18: data <= 32'hEA43AF00;	14'h2C19: data <= 32'hEA422890;	14'h2C1A: data <= 32'hEA40A221;	14'h2C1B: data <= 32'hEA3F1BB1;	14'h2C1C: data <= 32'hEA3D9541;	14'h2C1D: data <= 32'hEA3C0ED2;	14'h2C1E: data <= 32'hEA3A8862;	14'h2C1F: data <= 32'hEA3901F2;	14'h2C20: data <= 32'hEA377B82;	14'h2C21: data <= 32'hEA35F513;	14'h2C22: data <= 32'hEA346EA3;	14'h2C23: data <= 32'hEA32E833;	14'h2C24: data <= 32'hEA3161C3;	14'h2C25: data <= 32'hEA2FDB54;	14'h2C26: data <= 32'hEA2E54E4;	14'h2C27: data <= 32'hEA2C4723;	14'h2C28: data <= 32'hEA28F98D;	14'h2C29: data <= 32'hEA25ABF7;	14'h2C2A: data <= 32'hEA225E60;	14'h2C2B: data <= 32'hEA1F10CA;	14'h2C2C: data <= 32'hEA1BC334;	14'h2C2D: data <= 32'hEA18759D;	14'h2C2E: data <= 32'hEA152807;	14'h2C2F: data <= 32'hEA11DA71;	14'h2C30: data <= 32'hEA0E8CDA;	14'h2C31: data <= 32'hEA0B3F44;	14'h2C32: data <= 32'hEA07F1AE;	14'h2C33: data <= 32'hEA04A417;	14'h2C34: data <= 32'hEA015681;	14'h2C35: data <= 32'hE9FE08EB;	14'h2C36: data <= 32'hE9FABB54;	14'h2C37: data <= 32'hE9F75D5C;	14'h2C38: data <= 32'hE9F345B9;	14'h2C39: data <= 32'hE9EF2E15;	14'h2C3A: data <= 32'hE9EB1672;	14'h2C3B: data <= 32'hE9E6FECE;	14'h2C3C: data <= 32'hE9E2E72B;	14'h2C3D: data <= 32'hE9DECF88;	14'h2C3E: data <= 32'hE9DAB7E4;	14'h2C3F: data <= 32'hE9D6A041;	14'h2C40: data <= 32'hE9D2889E;	14'h2C41: data <= 32'hE9CE70FA;	14'h2C42: data <= 32'hE9CA5957;	14'h2C43: data <= 32'hE9C641B4;	14'h2C44: data <= 32'hE9C22A10;	14'h2C45: data <= 32'hE9BE126D;	14'h2C46: data <= 32'hE9B9FAC9;	14'h2C47: data <= 32'hE9B5E326;	14'h2C48: data <= 32'hE9B45277;	14'h2C49: data <= 32'hE9B326DF;	14'h2C4A: data <= 32'hE9B1FB47;	14'h2C4B: data <= 32'hE9B0CFAE;	14'h2C4C: data <= 32'hE9AFA416;	14'h2C4D: data <= 32'hE9AE787D;	14'h2C4E: data <= 32'hE9AD4CE5;	14'h2C4F: data <= 32'hE9AC214C;	14'h2C50: data <= 32'hE9AAF5B4;	14'h2C51: data <= 32'hE9A9CA1C;	14'h2C52: data <= 32'hE9A89E83;	14'h2C53: data <= 32'hE9A772EB;	14'h2C54: data <= 32'hE9A64752;	14'h2C55: data <= 32'hE9A51BBA;	14'h2C56: data <= 32'hE9A3F021;	14'h2C57: data <= 32'hE9A2C489;	14'h2C58: data <= 32'hE9A2BED6;	14'h2C59: data <= 32'hE9A35854;	14'h2C5A: data <= 32'hE9A3F1D2;	14'h2C5B: data <= 32'hE9A48B51;	14'h2C5C: data <= 32'hE9A524CF;	14'h2C5D: data <= 32'hE9A5BE4D;	14'h2C5E: data <= 32'hE9A657CC;	14'h2C5F: data <= 32'hE9A6F14A;	14'h2C60: data <= 32'hE9A78AC8;	14'h2C61: data <= 32'hE9A82446;	14'h2C62: data <= 32'hE9A8BDC5;	14'h2C63: data <= 32'hE9A95743;	14'h2C64: data <= 32'hE9A9F0C1;	14'h2C65: data <= 32'hE9AA8A40;	14'h2C66: data <= 32'hE9AB23BE;	14'h2C67: data <= 32'hE9ABBD3C;	14'h2C68: data <= 32'hE9AC3D58;	14'h2C69: data <= 32'hE9AC9C24;	14'h2C6A: data <= 32'hE9ACFAEF;	14'h2C6B: data <= 32'hE9AD59BB;	14'h2C6C: data <= 32'hE9ADB886;	14'h2C6D: data <= 32'hE9AE1751;	14'h2C6E: data <= 32'hE9AE761D;	14'h2C6F: data <= 32'hE9AED4E8;	14'h2C70: data <= 32'hE9AF33B3;	14'h2C71: data <= 32'hE9AF927F;	14'h2C72: data <= 32'hE9AFF14A;	14'h2C73: data <= 32'hE9B05016;	14'h2C74: data <= 32'hE9B0AEE1;	14'h2C75: data <= 32'hE9B10DAC;	14'h2C76: data <= 32'hE9B16C78;	14'h2C77: data <= 32'hE9B1CB43;	14'h2C78: data <= 32'hE9B219D6;	14'h2C79: data <= 32'hE9B22D9A;	14'h2C7A: data <= 32'hE9B2415E;	14'h2C7B: data <= 32'hE9B25523;	14'h2C7C: data <= 32'hE9B268E7;	14'h2C7D: data <= 32'hE9B27CAB;	14'h2C7E: data <= 32'hE9B2906F;	14'h2C7F: data <= 32'hE9B2A434;	14'h2C80: data <= 32'hE9B2B7F8;	14'h2C81: data <= 32'hE9B2CBBC;	14'h2C82: data <= 32'hE9B2DF81;	14'h2C83: data <= 32'hE9B2F345;	14'h2C84: data <= 32'hE9B30709;	14'h2C85: data <= 32'hE9B31ACE;	14'h2C86: data <= 32'hE9B32E92;	14'h2C87: data <= 32'hE9B34256;	14'h2C88: data <= 32'hE9B3561A;	14'h2C89: data <= 32'hE9B2A686;	14'h2C8A: data <= 32'hE9B1F6F1;	14'h2C8B: data <= 32'hE9B1475D;	14'h2C8C: data <= 32'hE9B097C8;	14'h2C8D: data <= 32'hE9AFE834;	14'h2C8E: data <= 32'hE9AF389F;	14'h2C8F: data <= 32'hE9AE890A;	14'h2C90: data <= 32'hE9ADD976;	14'h2C91: data <= 32'hE9AD29E1;	14'h2C92: data <= 32'hE9AC7A4D;	14'h2C93: data <= 32'hE9ABCAB8;	14'h2C94: data <= 32'hE9AB1B23;	14'h2C95: data <= 32'hE9AA6B8F;	14'h2C96: data <= 32'hE9A9BBFA;	14'h2C97: data <= 32'hE9A90C66;	14'h2C98: data <= 32'hE9A85CD1;	14'h2C99: data <= 32'hE9A80791;	14'h2C9A: data <= 32'hE9A7CB3C;	14'h2C9B: data <= 32'hE9A78EE7;	14'h2C9C: data <= 32'hE9A75292;	14'h2C9D: data <= 32'hE9A7163D;	14'h2C9E: data <= 32'hE9A6D9E8;	14'h2C9F: data <= 32'hE9A69D94;	14'h2CA0: data <= 32'hE9A6613F;	14'h2CA1: data <= 32'hE9A624EA;	14'h2CA2: data <= 32'hE9A5E895;	14'h2CA3: data <= 32'hE9A5AC40;	14'h2CA4: data <= 32'hE9A56FEB;	14'h2CA5: data <= 32'hE9A53396;	14'h2CA6: data <= 32'hE9A4F741;	14'h2CA7: data <= 32'hE9A4BAEC;	14'h2CA8: data <= 32'hE9A47E97;	14'h2CA9: data <= 32'hE9A36EF4;	14'h2CAA: data <= 32'hE9A1BE52;	14'h2CAB: data <= 32'hE9A00DAF;	14'h2CAC: data <= 32'hE99E5D0D;	14'h2CAD: data <= 32'hE99CAC6B;	14'h2CAE: data <= 32'hE99AFBC8;	14'h2CAF: data <= 32'hE9994B26;	14'h2CB0: data <= 32'hE9979A84;	14'h2CB1: data <= 32'hE995E9E1;	14'h2CB2: data <= 32'hE994393F;	14'h2CB3: data <= 32'hE992889D;	14'h2CB4: data <= 32'hE990D7FA;	14'h2CB5: data <= 32'hE98F2758;	14'h2CB6: data <= 32'hE98D76B6;	14'h2CB7: data <= 32'hE98BC613;	14'h2CB8: data <= 32'hE98A1571;	14'h2CB9: data <= 32'hE985CB52;	14'h2CBA: data <= 32'hE97CB499;	14'h2CBB: data <= 32'hE9739DE1;	14'h2CBC: data <= 32'hE96A8729;	14'h2CBD: data <= 32'hE9617071;	14'h2CBE: data <= 32'hE95859B9;	14'h2CBF: data <= 32'hE94F4301;	14'h2CC0: data <= 32'hE9462C49;	14'h2CC1: data <= 32'hE93D1591;	14'h2CC2: data <= 32'hE933FED8;	14'h2CC3: data <= 32'hE92AE820;	14'h2CC4: data <= 32'hE921D168;	14'h2CC5: data <= 32'hE918BAB0;	14'h2CC6: data <= 32'hE90FA3F8;	14'h2CC7: data <= 32'hE9068D40;	14'h2CC8: data <= 32'hE8FD7688;	14'h2CC9: data <= 32'hE8F3713D;	14'h2CCA: data <= 32'hE8E37517;	14'h2CCB: data <= 32'hE8D378F1;	14'h2CCC: data <= 32'hE8C37CCB;	14'h2CCD: data <= 32'hE8B380A5;	14'h2CCE: data <= 32'hE8A3847F;	14'h2CCF: data <= 32'hE8938859;	14'h2CD0: data <= 32'hE8838C33;	14'h2CD1: data <= 32'hE873900D;	14'h2CD2: data <= 32'hE86393E7;	14'h2CD3: data <= 32'hE85397C1;	14'h2CD4: data <= 32'hE8439B9B;	14'h2CD5: data <= 32'hE8339F75;	14'h2CD6: data <= 32'hE823A34F;	14'h2CD7: data <= 32'hE813A729;	14'h2CD8: data <= 32'hE803AB03;	14'h2CD9: data <= 32'hE7F3AEDD;	14'h2CDA: data <= 32'hE7E4ACFC;	14'h2CDB: data <= 32'hE7D5C130;	14'h2CDC: data <= 32'hE7C6D564;	14'h2CDD: data <= 32'hE7B7E998;	14'h2CDE: data <= 32'hE7A8FDCC;	14'h2CDF: data <= 32'hE79A1200;	14'h2CE0: data <= 32'hE78B2634;	14'h2CE1: data <= 32'hE77C3A68;	14'h2CE2: data <= 32'hE76D4E9C;	14'h2CE3: data <= 32'hE75E62D0;	14'h2CE4: data <= 32'hE74F7704;	14'h2CE5: data <= 32'hE7408B38;	14'h2CE6: data <= 32'hE7319F6C;	14'h2CE7: data <= 32'hE722B3A0;	14'h2CE8: data <= 32'hE713C7D4;	14'h2CE9: data <= 32'hE704DC08;	14'h2CEA: data <= 32'hE6F5B579;	14'h2CEB: data <= 32'hE6E6760E;	14'h2CEC: data <= 32'hE6D736A3;	14'h2CED: data <= 32'hE6C7F737;	14'h2CEE: data <= 32'hE6B8B7CC;	14'h2CEF: data <= 32'hE6A97861;	14'h2CF0: data <= 32'hE69A38F6;	14'h2CF1: data <= 32'hE68AF98B;	14'h2CF2: data <= 32'hE67BBA1F;	14'h2CF3: data <= 32'hE66C7AB4;	14'h2CF4: data <= 32'hE65D3B49;	14'h2CF5: data <= 32'hE64DFBDE;	14'h2CF6: data <= 32'hE63EBC72;	14'h2CF7: data <= 32'hE62F7D07;	14'h2CF8: data <= 32'hE6203D9C;	14'h2CF9: data <= 32'hE610FE31;	14'h2CFA: data <= 32'hE605215D;	14'h2CFB: data <= 32'hE5FCD746;	14'h2CFC: data <= 32'hE5F48D2F;	14'h2CFD: data <= 32'hE5EC4318;	14'h2CFE: data <= 32'hE5E3F901;	14'h2CFF: data <= 32'hE5DBAEEA;	14'h2D00: data <= 32'hE5D364D3;	14'h2D01: data <= 32'hE5CB1ABC;	14'h2D02: data <= 32'hE5C2D0A5;	14'h2D03: data <= 32'hE5BA868D;	14'h2D04: data <= 32'hE5B23C76;	14'h2D05: data <= 32'hE5A9F25F;	14'h2D06: data <= 32'hE5A1A848;	14'h2D07: data <= 32'hE5995E31;	14'h2D08: data <= 32'hE591141A;	14'h2D09: data <= 32'hE588CA03;	14'h2D0A: data <= 32'hE5838A89;	14'h2D0B: data <= 32'hE5868152;	14'h2D0C: data <= 32'hE589781B;	14'h2D0D: data <= 32'hE58C6EE4;	14'h2D0E: data <= 32'hE58F65AE;	14'h2D0F: data <= 32'hE5925C77;	14'h2D10: data <= 32'hE5955340;	14'h2D11: data <= 32'hE5984A09;	14'h2D12: data <= 32'hE59B40D2;	14'h2D13: data <= 32'hE59E379B;	14'h2D14: data <= 32'hE5A12E64;	14'h2D15: data <= 32'hE5A4252D;	14'h2D16: data <= 32'hE5A71BF6;	14'h2D17: data <= 32'hE5AA12BF;	14'h2D18: data <= 32'hE5AD0988;	14'h2D19: data <= 32'hE5B00051;	14'h2D1A: data <= 32'hE5B2E4CD;	14'h2D1B: data <= 32'hE5B488F9;	14'h2D1C: data <= 32'hE5B62D25;	14'h2D1D: data <= 32'hE5B7D151;	14'h2D1E: data <= 32'hE5B9757D;	14'h2D1F: data <= 32'hE5BB19AA;	14'h2D20: data <= 32'hE5BCBDD6;	14'h2D21: data <= 32'hE5BE6202;	14'h2D22: data <= 32'hE5C0062E;	14'h2D23: data <= 32'hE5C1AA5A;	14'h2D24: data <= 32'hE5C34E87;	14'h2D25: data <= 32'hE5C4F2B3;	14'h2D26: data <= 32'hE5C696DF;	14'h2D27: data <= 32'hE5C83B0B;	14'h2D28: data <= 32'hE5C9DF37;	14'h2D29: data <= 32'hE5CB8363;	14'h2D2A: data <= 32'hE5CD2790;	14'h2D2B: data <= 32'hE5C8E467;	14'h2D2C: data <= 32'hE5C37CBB;	14'h2D2D: data <= 32'hE5BE150F;	14'h2D2E: data <= 32'hE5B8AD62;	14'h2D2F: data <= 32'hE5B345B6;	14'h2D30: data <= 32'hE5ADDE0A;	14'h2D31: data <= 32'hE5A8765E;	14'h2D32: data <= 32'hE5A30EB1;	14'h2D33: data <= 32'hE59DA705;	14'h2D34: data <= 32'hE5983F59;	14'h2D35: data <= 32'hE592D7AC;	14'h2D36: data <= 32'hE58D7000;	14'h2D37: data <= 32'hE5880854;	14'h2D38: data <= 32'hE582A0A7;	14'h2D39: data <= 32'hE57D38FB;	14'h2D3A: data <= 32'hE577D14F;	14'h2D3B: data <= 32'hE5728B8F;	14'h2D3C: data <= 32'hE56D5A76;	14'h2D3D: data <= 32'hE568295C;	14'h2D3E: data <= 32'hE562F843;	14'h2D3F: data <= 32'hE55DC729;	14'h2D40: data <= 32'hE5589610;	14'h2D41: data <= 32'hE55364F6;	14'h2D42: data <= 32'hE54E33DD;	14'h2D43: data <= 32'hE54902C3;	14'h2D44: data <= 32'hE543D1AA;	14'h2D45: data <= 32'hE53EA090;	14'h2D46: data <= 32'hE5396F77;	14'h2D47: data <= 32'hE5343E5D;	14'h2D48: data <= 32'hE52F0D44;	14'h2D49: data <= 32'hE529DC2A;	14'h2D4A: data <= 32'hE524AB11;	14'h2D4B: data <= 32'hE51FB025;	14'h2D4C: data <= 32'hE51B04B0;	14'h2D4D: data <= 32'hE516593A;	14'h2D4E: data <= 32'hE511ADC5;	14'h2D4F: data <= 32'hE50D024F;	14'h2D50: data <= 32'hE50856D9;	14'h2D51: data <= 32'hE503AB64;	14'h2D52: data <= 32'hE4FEFFEE;	14'h2D53: data <= 32'hE4FA5479;	14'h2D54: data <= 32'hE4F5A903;	14'h2D55: data <= 32'hE4F0FD8E;	14'h2D56: data <= 32'hE4EC5218;	14'h2D57: data <= 32'hE4E7A6A3;	14'h2D58: data <= 32'hE4E2FB2D;	14'h2D59: data <= 32'hE4DE4FB8;	14'h2D5A: data <= 32'hE4D9A442;	14'h2D5B: data <= 32'hE4D3FDBD;	14'h2D5C: data <= 32'hE4CA233E;	14'h2D5D: data <= 32'hE4C048BF;	14'h2D5E: data <= 32'hE4B66E40;	14'h2D5F: data <= 32'hE4AC93C1;	14'h2D60: data <= 32'hE4A2B942;	14'h2D61: data <= 32'hE498DEC3;	14'h2D62: data <= 32'hE48F0444;	14'h2D63: data <= 32'hE48529C5;	14'h2D64: data <= 32'hE47B4F46;	14'h2D65: data <= 32'hE47174C7;	14'h2D66: data <= 32'hE4679A48;	14'h2D67: data <= 32'hE45DBFC9;	14'h2D68: data <= 32'hE453E54A;	14'h2D69: data <= 32'hE44A0ACB;	14'h2D6A: data <= 32'hE440304C;	14'h2D6B: data <= 32'hE43655CD;	14'h2D6C: data <= 32'hE42B4191;	14'h2D6D: data <= 32'hE420249D;	14'h2D6E: data <= 32'hE41507A9;	14'h2D6F: data <= 32'hE409EAB6;	14'h2D70: data <= 32'hE3FECDC2;	14'h2D71: data <= 32'hE3F3B0CE;	14'h2D72: data <= 32'hE3E893DB;	14'h2D73: data <= 32'hE3DD76E7;	14'h2D74: data <= 32'hE3D259F3;	14'h2D75: data <= 32'hE3C73D00;	14'h2D76: data <= 32'hE3BC200C;	14'h2D77: data <= 32'hE3B10318;	14'h2D78: data <= 32'hE3A5E624;	14'h2D79: data <= 32'hE39AC931;	14'h2D7A: data <= 32'hE38FAC3D;	14'h2D7B: data <= 32'hE3848F49;	14'h2D7C: data <= 32'hE37D6888;	14'h2D7D: data <= 32'hE37787C4;	14'h2D7E: data <= 32'hE371A6FF;	14'h2D7F: data <= 32'hE36BC63B;	14'h2D80: data <= 32'hE365E577;	14'h2D81: data <= 32'hE36004B3;	14'h2D82: data <= 32'hE35A23EF;	14'h2D83: data <= 32'hE354432B;	14'h2D84: data <= 32'hE34E6267;	14'h2D85: data <= 32'hE34881A3;	14'h2D86: data <= 32'hE342A0DF;	14'h2D87: data <= 32'hE33CC01B;	14'h2D88: data <= 32'hE336DF57;	14'h2D89: data <= 32'hE330FE93;	14'h2D8A: data <= 32'hE32B1DCF;	14'h2D8B: data <= 32'hE3253D0B;	14'h2D8C: data <= 32'hE322D4D4;	14'h2D8D: data <= 32'hE3235FE2;	14'h2D8E: data <= 32'hE323EAF0;	14'h2D8F: data <= 32'hE32475FE;	14'h2D90: data <= 32'hE325010C;	14'h2D91: data <= 32'hE3258C1A;	14'h2D92: data <= 32'hE3261728;	14'h2D93: data <= 32'hE326A236;	14'h2D94: data <= 32'hE3272D44;	14'h2D95: data <= 32'hE327B852;	14'h2D96: data <= 32'hE3284360;	14'h2D97: data <= 32'hE328CE6E;	14'h2D98: data <= 32'hE329597C;	14'h2D99: data <= 32'hE329E48A;	14'h2D9A: data <= 32'hE32A6F98;	14'h2D9B: data <= 32'hE32AFAA6;	14'h2D9C: data <= 32'hE32B0E4B;	14'h2D9D: data <= 32'hE32A292C;	14'h2D9E: data <= 32'hE329440C;	14'h2D9F: data <= 32'hE3285EED;	14'h2DA0: data <= 32'hE32779CE;	14'h2DA1: data <= 32'hE32694AE;	14'h2DA2: data <= 32'hE325AF8F;	14'h2DA3: data <= 32'hE324CA70;	14'h2DA4: data <= 32'hE323E550;	14'h2DA5: data <= 32'hE3230031;	14'h2DA6: data <= 32'hE3221B12;	14'h2DA7: data <= 32'hE32135F2;	14'h2DA8: data <= 32'hE32050D3;	14'h2DA9: data <= 32'hE31F6BB3;	14'h2DAA: data <= 32'hE31E8694;	14'h2DAB: data <= 32'hE31DA175;	14'h2DAC: data <= 32'hE31BB8E4;	14'h2DAD: data <= 32'hE31173E9;	14'h2DAE: data <= 32'hE3072EEF;	14'h2DAF: data <= 32'hE2FCE9F4;	14'h2DB0: data <= 32'hE2F2A4FA;	14'h2DB1: data <= 32'hE2E85FFF;	14'h2DB2: data <= 32'hE2DE1B05;	14'h2DB3: data <= 32'hE2D3D60A;	14'h2DB4: data <= 32'hE2C9910F;	14'h2DB5: data <= 32'hE2BF4C15;	14'h2DB6: data <= 32'hE2B5071A;	14'h2DB7: data <= 32'hE2AAC220;	14'h2DB8: data <= 32'hE2A07D25;	14'h2DB9: data <= 32'hE296382B;	14'h2DBA: data <= 32'hE28BF330;	14'h2DBB: data <= 32'hE281AE36;	14'h2DBC: data <= 32'hE277693B;	14'h2DBD: data <= 32'hE266EF0A;	14'h2DBE: data <= 32'hE255B438;	14'h2DBF: data <= 32'hE2447965;	14'h2DC0: data <= 32'hE2333E92;	14'h2DC1: data <= 32'hE22203C0;	14'h2DC2: data <= 32'hE210C8ED;	14'h2DC3: data <= 32'hE1FF8E1A;	14'h2DC4: data <= 32'hE1EE5348;	14'h2DC5: data <= 32'hE1DD1875;	14'h2DC6: data <= 32'hE1CBDDA2;	14'h2DC7: data <= 32'hE1BAA2CF;	14'h2DC8: data <= 32'hE1A967FD;	14'h2DC9: data <= 32'hE1982D2A;	14'h2DCA: data <= 32'hE186F257;	14'h2DCB: data <= 32'hE175B785;	14'h2DCC: data <= 32'hE1647CB2;	14'h2DCD: data <= 32'hE1504E29;	14'h2DCE: data <= 32'hE13AB4E2;	14'h2DCF: data <= 32'hE1251B9B;	14'h2DD0: data <= 32'hE10F8254;	14'h2DD1: data <= 32'hE0F9E90D;	14'h2DD2: data <= 32'hE0E44FC6;	14'h2DD3: data <= 32'hE0CEB67F;	14'h2DD4: data <= 32'hE0B91D37;	14'h2DD5: data <= 32'hE0A383F0;	14'h2DD6: data <= 32'hE08DEAA9;	14'h2DD7: data <= 32'hE0785162;	14'h2DD8: data <= 32'hE062B81B;	14'h2DD9: data <= 32'hE04D1ED4;	14'h2DDA: data <= 32'hE037858D;	14'h2DDB: data <= 32'hE021EC46;	14'h2DDC: data <= 32'hE00C52FF;	14'h2DDD: data <= 32'hDFF5FC61;	14'h2DDE: data <= 32'hDFDEC702;	14'h2DDF: data <= 32'hDFC791A3;	14'h2DE0: data <= 32'hDFB05C44;	14'h2DE1: data <= 32'hDF9926E4;	14'h2DE2: data <= 32'hDF81F185;	14'h2DE3: data <= 32'hDF6ABC26;	14'h2DE4: data <= 32'hDF5386C7;	14'h2DE5: data <= 32'hDF3C5168;	14'h2DE6: data <= 32'hDF251C09;	14'h2DE7: data <= 32'hDF0DE6AA;	14'h2DE8: data <= 32'hDEF6B14B;	14'h2DE9: data <= 32'hDEDF7BEC;	14'h2DEA: data <= 32'hDEC8468D;	14'h2DEB: data <= 32'hDEB1112E;	14'h2DEC: data <= 32'hDE99DBCF;	14'h2DED: data <= 32'hDE833B5D;	14'h2DEE: data <= 32'hDE6E6A3F;	14'h2DEF: data <= 32'hDE599921;	14'h2DF0: data <= 32'hDE44C803;	14'h2DF1: data <= 32'hDE2FF6E4;	14'h2DF2: data <= 32'hDE1B25C6;	14'h2DF3: data <= 32'hDE0654A8;	14'h2DF4: data <= 32'hDDF1838A;	14'h2DF5: data <= 32'hDDDCB26C;	14'h2DF6: data <= 32'hDDC7E14E;	14'h2DF7: data <= 32'hDDB31030;	14'h2DF8: data <= 32'hDD9E3F11;	14'h2DF9: data <= 32'hDD896DF3;	14'h2DFA: data <= 32'hDD749CD5;	14'h2DFB: data <= 32'hDD5FCBB7;	14'h2DFC: data <= 32'hDD4AFA99;	14'h2DFD: data <= 32'hDD360820;	14'h2DFE: data <= 32'hDD1C64F6;	14'h2DFF: data <= 32'hDD02C1CC;	14'h2E00: data <= 32'hDCE91EA2;	14'h2E01: data <= 32'hDCCF7B78;	14'h2E02: data <= 32'hDCB5D84D;	14'h2E03: data <= 32'hDC9C3523;	14'h2E04: data <= 32'hDC8291F9;	14'h2E05: data <= 32'hDC68EECF;	14'h2E06: data <= 32'hDC4F4BA4;	14'h2E07: data <= 32'hDC35A87A;	14'h2E08: data <= 32'hDC1C0550;	14'h2E09: data <= 32'hDC026226;	14'h2E0A: data <= 32'hDBE8BEFB;	14'h2E0B: data <= 32'hDBCF1BD1;	14'h2E0C: data <= 32'hDBB578A7;	14'h2E0D: data <= 32'hDB9BD57D;	14'h2E0E: data <= 32'hDB749749;	14'h2E0F: data <= 32'hDB4A2C60;	14'h2E10: data <= 32'hDB1FC176;	14'h2E11: data <= 32'hDAF5568D;	14'h2E12: data <= 32'hDACAEBA4;	14'h2E13: data <= 32'hDAA080BB;	14'h2E14: data <= 32'hDA7615D1;	14'h2E15: data <= 32'hDA4BAAE8;	14'h2E16: data <= 32'hDA213FFF;	14'h2E17: data <= 32'hD9F6D516;	14'h2E18: data <= 32'hD9CC6A2D;	14'h2E19: data <= 32'hD9A1FF43;	14'h2E1A: data <= 32'hD977945A;	14'h2E1B: data <= 32'hD94D2971;	14'h2E1C: data <= 32'hD922BE88;	14'h2E1D: data <= 32'hD8F8539E;	14'h2E1E: data <= 32'hD8C66E1C;	14'h2E1F: data <= 32'hD88F6F32;	14'h2E20: data <= 32'hD8587048;	14'h2E21: data <= 32'hD821715D;	14'h2E22: data <= 32'hD7EA7273;	14'h2E23: data <= 32'hD7B37388;	14'h2E24: data <= 32'hD77C749E;	14'h2E25: data <= 32'hD74575B4;	14'h2E26: data <= 32'hD70E76C9;	14'h2E27: data <= 32'hD6D777DF;	14'h2E28: data <= 32'hD6A078F4;	14'h2E29: data <= 32'hD6697A0A;	14'h2E2A: data <= 32'hD6327B20;	14'h2E2B: data <= 32'hD5FB7C35;	14'h2E2C: data <= 32'hD5C47D4B;	14'h2E2D: data <= 32'hD58D7E61;	14'h2E2E: data <= 32'hD555C747;	14'h2E2F: data <= 32'hD51CE195;	14'h2E30: data <= 32'hD4E3FBE3;	14'h2E31: data <= 32'hD4AB1632;	14'h2E32: data <= 32'hD4723080;	14'h2E33: data <= 32'hD4394ACF;	14'h2E34: data <= 32'hD400651D;	14'h2E35: data <= 32'hD3C77F6C;	14'h2E36: data <= 32'hD38E99BA;	14'h2E37: data <= 32'hD355B408;	14'h2E38: data <= 32'hD31CCE57;	14'h2E39: data <= 32'hD2E3E8A5;	14'h2E3A: data <= 32'hD2AB02F4;	14'h2E3B: data <= 32'hD2721D42;	14'h2E3C: data <= 32'hD2393791;	14'h2E3D: data <= 32'hD20051DF;	14'h2E3E: data <= 32'hD1CBE98B;	14'h2E3F: data <= 32'hD1AEB39B;	14'h2E40: data <= 32'hD1917DAC;	14'h2E41: data <= 32'hD17447BC;	14'h2E42: data <= 32'hD15711CD;	14'h2E43: data <= 32'hD139DBDD;	14'h2E44: data <= 32'hD11CA5ED;	14'h2E45: data <= 32'hD0FF6FFE;	14'h2E46: data <= 32'hD0E23A0E;	14'h2E47: data <= 32'hD0C5041E;	14'h2E48: data <= 32'hD0A7CE2F;	14'h2E49: data <= 32'hD08A983F;	14'h2E4A: data <= 32'hD06D624F;	14'h2E4B: data <= 32'hD0502C60;	14'h2E4C: data <= 32'hD032F670;	14'h2E4D: data <= 32'hD015C081;	14'h2E4E: data <= 32'hCFF88A91;	14'h2E4F: data <= 32'hCFEC1464;	14'h2E50: data <= 32'hCFE0933B;	14'h2E51: data <= 32'hCFD51212;	14'h2E52: data <= 32'hCFC990E9;	14'h2E53: data <= 32'hCFBE0FBF;	14'h2E54: data <= 32'hCFB28E96;	14'h2E55: data <= 32'hCFA70D6D;	14'h2E56: data <= 32'hCF9B8C44;	14'h2E57: data <= 32'hCF900B1B;	14'h2E58: data <= 32'hCF8489F2;	14'h2E59: data <= 32'hCF7908C9;	14'h2E5A: data <= 32'hCF6D879F;	14'h2E5B: data <= 32'hCF620676;	14'h2E5C: data <= 32'hCF56854D;	14'h2E5D: data <= 32'hCF4B0424;	14'h2E5E: data <= 32'hCF3F82FB;	14'h2E5F: data <= 32'hCF2A3016;	14'h2E60: data <= 32'hCF113A2E;	14'h2E61: data <= 32'hCEF84447;	14'h2E62: data <= 32'hCEDF4E5F;	14'h2E63: data <= 32'hCEC65877;	14'h2E64: data <= 32'hCEAD6290;	14'h2E65: data <= 32'hCE946CA8;	14'h2E66: data <= 32'hCE7B76C0;	14'h2E67: data <= 32'hCE6280D9;	14'h2E68: data <= 32'hCE498AF1;	14'h2E69: data <= 32'hCE309509;	14'h2E6A: data <= 32'hCE179F22;	14'h2E6B: data <= 32'hCDFEA93A;	14'h2E6C: data <= 32'hCDE5B352;	14'h2E6D: data <= 32'hCDCCBD6A;	14'h2E6E: data <= 32'hCDB3C783;	14'h2E6F: data <= 32'hCD9973B9;	14'h2E70: data <= 32'hCD7DD477;	14'h2E71: data <= 32'hCD623535;	14'h2E72: data <= 32'hCD4695F4;	14'h2E73: data <= 32'hCD2AF6B2;	14'h2E74: data <= 32'hCD0F5770;	14'h2E75: data <= 32'hCCF3B82F;	14'h2E76: data <= 32'hCCD818ED;	14'h2E77: data <= 32'hCCBC79AB;	14'h2E78: data <= 32'hCCA0DA6A;	14'h2E79: data <= 32'hCC853B28;	14'h2E7A: data <= 32'hCC699BE6;	14'h2E7B: data <= 32'hCC4DFCA4;	14'h2E7C: data <= 32'hCC325D63;	14'h2E7D: data <= 32'hCC16BE21;	14'h2E7E: data <= 32'hCBFB1EDF;	14'h2E7F: data <= 32'hCBDC275E;	14'h2E80: data <= 32'hCBB54803;	14'h2E81: data <= 32'hCB8E68A7;	14'h2E82: data <= 32'hCB67894B;	14'h2E83: data <= 32'hCB40A9EF;	14'h2E84: data <= 32'hCB19CA93;	14'h2E85: data <= 32'hCAF2EB37;	14'h2E86: data <= 32'hCACC0BDB;	14'h2E87: data <= 32'hCAA52C7F;	14'h2E88: data <= 32'hCA7E4D24;	14'h2E89: data <= 32'hCA576DC8;	14'h2E8A: data <= 32'hCA308E6C;	14'h2E8B: data <= 32'hCA09AF10;	14'h2E8C: data <= 32'hC9E2CFB4;	14'h2E8D: data <= 32'hC9BBF058;	14'h2E8E: data <= 32'hC99510FC;	14'h2E8F: data <= 32'hC96DB81A;	14'h2E90: data <= 32'hC940FDE8;	14'h2E91: data <= 32'hC91443B6;	14'h2E92: data <= 32'hC8E78984;	14'h2E93: data <= 32'hC8BACF52;	14'h2E94: data <= 32'hC88E1520;	14'h2E95: data <= 32'hC8615AEE;	14'h2E96: data <= 32'hC834A0BC;	14'h2E97: data <= 32'hC807E68A;	14'h2E98: data <= 32'hC7DB2C59;	14'h2E99: data <= 32'hC7AE7227;	14'h2E9A: data <= 32'hC781B7F5;	14'h2E9B: data <= 32'hC754FDC3;	14'h2E9C: data <= 32'hC7284391;	14'h2E9D: data <= 32'hC6FB895F;	14'h2E9E: data <= 32'hC6CECF2D;	14'h2E9F: data <= 32'hC6A214FB;	14'h2EA0: data <= 32'hC6666BD8;	14'h2EA1: data <= 32'hC6286D60;	14'h2EA2: data <= 32'hC5EA6EE7;	14'h2EA3: data <= 32'hC5AC706E;	14'h2EA4: data <= 32'hC56E71F6;	14'h2EA5: data <= 32'hC530737D;	14'h2EA6: data <= 32'hC4F27504;	14'h2EA7: data <= 32'hC4B4768C;	14'h2EA8: data <= 32'hC4767813;	14'h2EA9: data <= 32'hC438799A;	14'h2EAA: data <= 32'hC3FA7B21;	14'h2EAB: data <= 32'hC3BC7CA9;	14'h2EAC: data <= 32'hC37E7E30;	14'h2EAD: data <= 32'hC3407FB7;	14'h2EAE: data <= 32'hC302813F;	14'h2EAF: data <= 32'hC2C482C6;	14'h2EB0: data <= 32'hC264273C;	14'h2EB1: data <= 32'hC1F12E9F;	14'h2EB2: data <= 32'hC17E3601;	14'h2EB3: data <= 32'hC10B3D64;	14'h2EB4: data <= 32'hC09844C6;	14'h2EB5: data <= 32'hC0254C29;	14'h2EB6: data <= 32'hBFB2538B;	14'h2EB7: data <= 32'hBF3F5AEE;	14'h2EB8: data <= 32'hBECC6250;	14'h2EB9: data <= 32'hBE5969B3;	14'h2EBA: data <= 32'hBDE67115;	14'h2EBB: data <= 32'hBD737878;	14'h2EBC: data <= 32'hBD007FDA;	14'h2EBD: data <= 32'hBC8D873D;	14'h2EBE: data <= 32'hBC1A8E9F;	14'h2EBF: data <= 32'hBBA79602;	14'h2EC0: data <= 32'hBAF8E96E;	14'h2EC1: data <= 32'hB9FBE0A6;	14'h2EC2: data <= 32'hB8FED7DE;	14'h2EC3: data <= 32'hB801CF17;	14'h2EC4: data <= 32'hB704C64F;	14'h2EC5: data <= 32'hB607BD87;	14'h2EC6: data <= 32'hB50AB4BF;	14'h2EC7: data <= 32'hB40DABF8;	14'h2EC8: data <= 32'hB310A330;	14'h2EC9: data <= 32'hB2139A68;	14'h2ECA: data <= 32'hB11691A1;	14'h2ECB: data <= 32'hB01988D9;	14'h2ECC: data <= 32'hAF1C8011;	14'h2ECD: data <= 32'hAE1F7749;	14'h2ECE: data <= 32'hAD226E82;	14'h2ECF: data <= 32'hAC2565BA;	14'h2ED0: data <= 32'hAAEE7F2B;	14'h2ED1: data <= 32'hA8E5D4A9;	14'h2ED2: data <= 32'hA6DD2A26;	14'h2ED3: data <= 32'hA4D47FA4;	14'h2ED4: data <= 32'hA2CBD522;	14'h2ED5: data <= 32'hA0C32AA0;	14'h2ED6: data <= 32'h9EBA801E;	14'h2ED7: data <= 32'h9CB1D59B;	14'h2ED8: data <= 32'h9AA92B19;	14'h2ED9: data <= 32'h98A08097;	14'h2EDA: data <= 32'h9697D615;	14'h2EDB: data <= 32'h948F2B93;	14'h2EDC: data <= 32'h92868110;	14'h2EDD: data <= 32'h907DD68E;	14'h2EDE: data <= 32'h8E752C0C;	14'h2EDF: data <= 32'h8C6C818A; default: data <= 32'h0; endcase
    end
    endmodule